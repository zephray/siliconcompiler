# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# Standard density, single height
SITE unit
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.48 BY 3.33 ;
END unit

# Standard density, double height
SITE unitdbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.48 BY 6.66 ;
END unitdbl

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.48 ;
  MINWIDTH 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  EDGECAPACITANCE 40.697E-6 ;
  CAPACITANCE CPERSQDIST 36.9866E-6 ;
  RESISTANCE RPERSQ 12.8 ;

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5
  RESISTANCE 9.30 ;

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.37 ;
  MINENCLOSEDAREA 0.14 ;
  MINWIDTH 0.14 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 40.567E-6 ;
  CAPACITANCE CPERSQDIST 25.7784E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5
  RESISTANCE 9.00 ;

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.48 ;
  MINENCLOSEDAREA 0.14 ;
  MINWIDTH 0.14 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;

  EDGECAPACITANCE 32.918E-6 ;
  CAPACITANCE CPERSQDIST 14.7703E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  RESISTANCE 3.41 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.74 ;
  MINWIDTH 0.3 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 37.065E-6 ;
  CAPACITANCE CPERSQDIST 11.1883E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  RESISTANCE 3.41 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.96 ;
  MINWIDTH 0.3 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 34.169E-6 ;
  CAPACITANCE CPERSQDIST 7.84019E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  RESISTANCE 0.38 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.33 ;
  MINWIDTH 1.6 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 36.828E-6 ;
  CAPACITANCE CPERSQDIST 5.99155E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###

MACRO sky130_fd_sc_hs__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2bb2o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.180 1.335 1.620 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.180 1.850 1.620 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.255 4.195 0.670 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.450 3.235 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.065 1.310 3.960 1.400 ;
        RECT 0.250 0.245 3.960 1.310 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.820 0.560 2.980 ;
        RECT 0.125 1.150 0.295 1.820 ;
        RECT 0.125 0.420 0.590 1.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.760 2.130 1.090 3.245 ;
        RECT 1.325 2.905 2.515 3.075 ;
        RECT 1.325 1.960 1.495 2.905 ;
        RECT 1.665 2.300 1.995 2.735 ;
        RECT 2.185 2.470 2.515 2.905 ;
        RECT 1.665 2.130 2.530 2.300 ;
        RECT 0.730 1.790 2.190 1.960 ;
        RECT 0.730 1.650 0.900 1.790 ;
        RECT 0.465 1.320 0.900 1.650 ;
        RECT 2.020 1.210 2.190 1.790 ;
        RECT 2.360 1.780 2.530 2.130 ;
        RECT 2.715 2.120 2.885 2.980 ;
        RECT 3.085 2.290 3.445 3.245 ;
        RECT 3.645 2.120 3.895 2.980 ;
        RECT 2.715 1.950 3.895 2.120 ;
        RECT 3.645 1.940 3.895 1.950 ;
        RECT 2.360 1.450 2.665 1.780 ;
        RECT 2.020 1.030 2.900 1.210 ;
        RECT 3.540 1.010 3.870 1.290 ;
        RECT 0.770 0.085 1.100 1.010 ;
        RECT 1.285 0.520 1.590 1.010 ;
        RECT 1.760 0.690 2.935 0.860 ;
        RECT 1.285 0.255 2.595 0.520 ;
        RECT 2.765 0.085 2.935 0.690 ;
        RECT 3.145 0.840 3.870 1.010 ;
        RECT 3.145 0.085 3.315 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a2bb2o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a2bb2o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2bb2o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.180 3.255 2.150 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.385 1.180 2.755 1.510 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.180 1.315 1.550 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.180 1.050 2.025 1.240 ;
        RECT 3.085 1.050 4.440 1.240 ;
        RECT 0.180 0.245 4.440 1.050 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.350 3.920 2.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.265 1.890 0.515 2.980 ;
        RECT 0.715 2.060 1.045 3.245 ;
        RECT 1.245 1.890 1.415 2.980 ;
        RECT 0.265 1.720 1.415 1.890 ;
        RECT 1.585 2.810 2.920 2.980 ;
        RECT 1.585 2.020 1.945 2.810 ;
        RECT 1.585 1.550 1.755 2.020 ;
        RECT 2.265 1.850 2.580 2.640 ;
        RECT 2.750 2.490 2.920 2.810 ;
        RECT 3.105 2.660 3.495 3.245 ;
        RECT 4.065 2.660 4.395 3.245 ;
        RECT 2.750 2.320 4.470 2.490 ;
        RECT 1.485 1.380 1.755 1.550 ;
        RECT 1.925 1.680 2.580 1.850 ;
        RECT 1.485 1.010 1.655 1.380 ;
        RECT 0.290 0.085 0.620 1.010 ;
        RECT 1.080 0.840 1.655 1.010 ;
        RECT 1.925 1.010 2.175 1.680 ;
        RECT 4.090 1.350 4.470 2.320 ;
        RECT 1.925 0.840 2.870 1.010 ;
        RECT 1.080 0.350 1.480 0.840 ;
        RECT 1.650 0.085 2.520 0.670 ;
        RECT 2.690 0.350 2.870 0.840 ;
        RECT 3.050 0.085 3.315 0.940 ;
        RECT 4.100 0.085 4.350 1.130 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__a2bb2o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2bb2o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.350 2.850 1.780 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 3.360 1.350 3.685 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.260 7.075 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.260 6.115 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.415 1.140 4.905 1.240 ;
        RECT 0.415 0.245 7.185 1.140 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 1.010 1.970 1.340 2.980 ;
        RECT 1.910 1.970 2.240 2.980 ;
        RECT 0.665 1.800 2.240 1.970 ;
        RECT 0.665 1.780 0.835 1.800 ;
        RECT 0.125 1.130 0.835 1.780 ;
        RECT 0.125 0.960 2.045 1.130 ;
        RECT 0.935 0.350 1.185 0.960 ;
        RECT 1.795 0.350 2.045 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.560 2.140 0.810 3.245 ;
        RECT 1.540 2.140 1.710 3.245 ;
        RECT 2.410 1.950 2.780 3.245 ;
        RECT 3.290 2.120 3.620 2.980 ;
        RECT 4.060 2.905 5.210 3.075 ;
        RECT 4.060 2.290 4.390 2.905 ;
        RECT 3.020 1.950 4.150 2.120 ;
        RECT 1.035 1.300 2.385 1.630 ;
        RECT 2.215 1.180 2.385 1.300 ;
        RECT 2.215 1.010 2.815 1.180 ;
        RECT 3.020 1.130 3.190 1.950 ;
        RECT 3.855 1.470 4.150 1.950 ;
        RECT 4.565 1.180 4.760 2.735 ;
        RECT 4.960 2.120 5.210 2.905 ;
        RECT 5.410 2.290 5.660 3.245 ;
        RECT 5.860 2.120 6.190 2.980 ;
        RECT 6.390 2.290 6.560 3.245 ;
        RECT 6.760 2.120 7.090 2.980 ;
        RECT 4.960 1.950 7.090 2.120 ;
        RECT 0.505 0.085 0.755 0.790 ;
        RECT 1.365 0.085 1.615 0.790 ;
        RECT 2.225 0.085 2.475 0.840 ;
        RECT 2.645 0.425 2.815 1.010 ;
        RECT 2.985 0.595 3.190 1.130 ;
        RECT 3.360 1.010 4.815 1.180 ;
        RECT 3.360 0.425 3.530 1.010 ;
        RECT 2.645 0.255 3.530 0.425 ;
        RECT 3.700 0.085 4.385 0.840 ;
        RECT 4.565 0.600 4.815 1.010 ;
        RECT 5.005 0.920 7.095 1.090 ;
        RECT 5.005 0.770 6.115 0.920 ;
        RECT 4.565 0.350 5.765 0.600 ;
        RECT 5.945 0.350 6.115 0.770 ;
        RECT 6.295 0.350 6.665 0.750 ;
        RECT 6.845 0.350 7.095 0.920 ;
        RECT 6.495 0.085 6.665 0.350 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__a2bb2o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2bb2oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.260 0.435 1.780 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.450 1.100 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.180 3.255 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.540 2.755 2.150 ;
        RECT 2.220 1.220 2.755 1.540 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.085 0.245 3.305 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.515200 ;
    PORT
      LAYER li1 ;
        RECT 1.530 2.290 1.780 2.980 ;
        RECT 1.610 2.220 1.780 2.290 ;
        RECT 1.610 1.920 2.275 2.220 ;
        RECT 1.610 1.750 2.050 1.920 ;
        RECT 1.880 1.050 2.050 1.750 ;
        RECT 1.880 0.880 2.315 1.050 ;
        RECT 2.055 0.350 2.315 0.880 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.120 1.950 0.450 3.245 ;
        RECT 2.430 2.980 2.600 3.245 ;
        RECT 0.960 2.120 1.290 2.980 ;
        RECT 1.980 2.560 2.230 2.980 ;
        RECT 2.430 2.730 2.790 2.980 ;
        RECT 2.990 2.560 3.240 2.980 ;
        RECT 1.980 2.390 3.240 2.560 ;
        RECT 0.960 1.950 1.440 2.120 ;
        RECT 1.270 1.550 1.440 1.950 ;
        RECT 2.990 1.820 3.240 2.390 ;
        RECT 1.270 1.220 1.710 1.550 ;
        RECT 1.270 1.130 1.440 1.220 ;
        RECT 0.175 0.085 0.425 1.090 ;
        RECT 0.605 0.960 1.440 1.130 ;
        RECT 0.605 0.540 0.935 0.960 ;
        RECT 1.105 0.710 1.710 0.790 ;
        RECT 1.105 0.085 1.885 0.710 ;
        RECT 2.885 0.085 3.215 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a2bb2oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a2bb2oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2bb2oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.285 0.435 0.670 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.450 1.570 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 4.675 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.320 3.735 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.515 1.240 2.850 1.280 ;
        RECT 0.515 0.245 5.175 1.240 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.750400 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.410 2.780 2.735 ;
        RECT 2.525 1.150 3.235 1.410 ;
        RECT 2.080 0.980 3.795 1.150 ;
        RECT 2.080 0.390 2.250 0.980 ;
        RECT 3.465 0.770 3.795 0.980 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.580 1.940 0.910 3.245 ;
        RECT 1.420 1.950 1.910 2.980 ;
        RECT 1.740 1.650 1.910 1.950 ;
        RECT 2.080 2.905 3.230 3.075 ;
        RECT 2.080 1.820 2.330 2.905 ;
        RECT 2.980 2.120 3.230 2.905 ;
        RECT 3.430 2.290 3.760 3.245 ;
        RECT 3.960 2.120 4.130 2.980 ;
        RECT 4.330 2.290 4.660 3.245 ;
        RECT 4.860 2.120 5.110 2.980 ;
        RECT 2.980 1.950 5.110 2.120 ;
        RECT 2.980 1.820 3.230 1.950 ;
        RECT 4.860 1.820 5.110 1.950 ;
        RECT 1.740 1.320 2.205 1.650 ;
        RECT 1.740 1.280 1.910 1.320 ;
        RECT 0.605 0.085 0.855 1.170 ;
        RECT 1.035 1.110 1.910 1.280 ;
        RECT 1.035 0.490 1.330 1.110 ;
        RECT 3.975 1.010 5.085 1.180 ;
        RECT 1.570 0.085 1.900 0.940 ;
        RECT 2.430 0.085 2.760 0.810 ;
        RECT 3.975 0.600 4.145 1.010 ;
        RECT 3.035 0.350 4.145 0.600 ;
        RECT 4.325 0.085 4.575 0.840 ;
        RECT 4.755 0.350 5.085 1.010 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__a2bb2oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2bb2oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.470 2.275 1.800 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.420 0.455 1.770 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.735 1.350 8.515 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 6.115 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.850 0.245 8.390 1.240 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.500800 ;
    PORT
      LAYER li1 ;
        RECT 3.185 1.890 3.355 2.735 ;
        RECT 4.085 1.890 4.255 2.735 ;
        RECT 3.185 1.720 4.255 1.890 ;
        RECT 3.965 1.130 4.255 1.720 ;
        RECT 3.965 0.960 6.150 1.130 ;
        RECT 2.270 0.790 6.150 0.960 ;
        RECT 2.270 0.350 2.520 0.790 ;
        RECT 3.210 0.350 3.380 0.790 ;
        RECT 4.960 0.770 6.150 0.790 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.105 2.905 1.255 3.075 ;
        RECT 0.105 1.940 0.435 2.905 ;
        RECT 0.635 1.300 0.885 2.735 ;
        RECT 1.085 2.140 1.255 2.905 ;
        RECT 1.455 2.310 1.705 3.245 ;
        RECT 1.905 2.140 2.235 2.980 ;
        RECT 1.085 1.970 2.235 2.140 ;
        RECT 2.655 2.905 4.785 3.075 ;
        RECT 1.085 1.940 1.255 1.970 ;
        RECT 2.655 1.820 2.985 2.905 ;
        RECT 3.555 2.060 3.885 2.905 ;
        RECT 4.455 2.120 4.785 2.905 ;
        RECT 4.985 2.290 5.155 3.245 ;
        RECT 5.355 2.120 5.685 2.980 ;
        RECT 5.885 2.290 6.135 3.245 ;
        RECT 6.335 2.120 6.505 2.980 ;
        RECT 6.705 2.290 6.955 3.245 ;
        RECT 7.155 2.120 7.485 2.980 ;
        RECT 7.685 2.290 7.855 3.245 ;
        RECT 8.055 2.120 8.385 2.980 ;
        RECT 4.455 1.950 8.385 2.120 ;
        RECT 6.335 1.820 6.505 1.950 ;
        RECT 2.575 1.300 3.585 1.550 ;
        RECT 0.635 1.130 3.585 1.300 ;
        RECT 0.940 0.085 1.270 0.960 ;
        RECT 1.450 0.350 1.620 1.130 ;
        RECT 6.330 1.010 8.300 1.180 ;
        RECT 1.800 0.085 2.090 0.885 ;
        RECT 2.700 0.085 3.030 0.620 ;
        RECT 3.560 0.085 3.890 0.620 ;
        RECT 6.330 0.600 6.500 1.010 ;
        RECT 4.530 0.350 6.500 0.600 ;
        RECT 6.680 0.085 6.930 0.840 ;
        RECT 7.110 0.350 7.360 1.010 ;
        RECT 7.540 0.085 7.790 0.840 ;
        RECT 7.970 0.350 8.300 1.010 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__a2bb2oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21bo_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.450 1.315 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 0.435 0.670 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.180 2.845 1.550 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.065 1.050 1.905 1.450 ;
        RECT 2.790 1.050 3.715 1.240 ;
        RECT 0.065 0.245 3.715 1.050 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 3.430 1.820 3.755 2.980 ;
        RECT 3.585 1.130 3.755 1.820 ;
        RECT 3.295 0.350 3.755 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.130 2.120 0.460 2.980 ;
        RECT 0.660 2.290 0.860 3.245 ;
        RECT 1.060 2.120 1.390 2.980 ;
        RECT 0.130 1.950 1.390 2.120 ;
        RECT 1.575 2.410 1.760 2.980 ;
        RECT 2.900 2.580 3.230 3.245 ;
        RECT 1.575 2.240 3.255 2.410 ;
        RECT 0.130 1.940 0.460 1.950 ;
        RECT 1.575 1.940 1.760 2.240 ;
        RECT 0.155 1.095 0.485 1.340 ;
        RECT 1.575 1.280 1.745 1.940 ;
        RECT 2.075 1.820 2.695 2.070 ;
        RECT 2.075 1.770 2.245 1.820 ;
        RECT 0.945 1.110 1.745 1.280 ;
        RECT 0.155 0.840 0.775 1.095 ;
        RECT 0.605 0.085 0.775 0.840 ;
        RECT 0.945 0.660 1.315 1.110 ;
        RECT 1.915 1.100 2.245 1.770 ;
        RECT 3.085 1.650 3.255 2.240 ;
        RECT 3.085 1.320 3.415 1.650 ;
        RECT 2.075 0.940 2.245 1.100 ;
        RECT 1.485 0.085 1.815 0.930 ;
        RECT 2.075 0.350 2.720 0.940 ;
        RECT 2.900 0.085 3.115 0.895 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a21bo_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21bo_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.725 1.260 3.235 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.450 3.735 1.780 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.510 1.550 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.180 0.245 3.820 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.020 1.820 1.415 2.070 ;
        RECT 1.020 1.040 1.190 1.820 ;
        RECT 1.020 0.840 1.395 1.040 ;
        RECT 1.225 0.750 1.395 0.840 ;
        RECT 1.225 0.350 1.565 0.750 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.120 2.410 0.450 2.700 ;
        RECT 0.635 2.580 0.965 3.245 ;
        RECT 1.535 2.580 1.865 3.245 ;
        RECT 0.120 2.240 1.810 2.410 ;
        RECT 0.120 1.820 0.450 2.240 ;
        RECT 0.680 1.010 0.850 2.240 ;
        RECT 1.605 1.890 1.810 2.240 ;
        RECT 2.055 2.060 2.415 2.980 ;
        RECT 2.585 2.270 2.755 2.980 ;
        RECT 2.955 2.440 3.205 3.245 ;
        RECT 3.405 2.270 3.735 2.980 ;
        RECT 2.585 2.100 3.735 2.270 ;
        RECT 2.245 1.930 2.415 2.060 ;
        RECT 3.405 1.950 3.735 2.100 ;
        RECT 1.605 1.720 2.075 1.890 ;
        RECT 2.245 1.760 2.555 1.930 ;
        RECT 1.905 1.590 2.075 1.720 ;
        RECT 1.360 1.220 1.735 1.550 ;
        RECT 1.905 1.260 2.215 1.590 ;
        RECT 0.270 0.840 0.850 1.010 ;
        RECT 1.565 1.090 1.735 1.220 ;
        RECT 2.385 1.090 2.555 1.760 ;
        RECT 1.565 0.920 2.810 1.090 ;
        RECT 0.270 0.540 0.600 0.840 ;
        RECT 0.805 0.085 1.055 0.670 ;
        RECT 1.735 0.085 2.310 0.750 ;
        RECT 2.480 0.350 2.810 0.920 ;
        RECT 3.380 0.085 3.710 1.090 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a21bo_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21bo_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.450 5.200 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.935 0.255 4.265 0.670 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.505 0.355 0.670 ;
        RECT 0.125 0.255 0.625 0.505 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.195 1.370 1.235 1.385 ;
        RECT 2.580 1.370 6.065 1.385 ;
        RECT 0.195 0.245 6.065 1.370 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.850 2.300 2.100 ;
        RECT 0.605 1.510 1.420 1.850 ;
        RECT 1.250 1.180 1.420 1.510 ;
        RECT 1.250 1.010 2.415 1.180 ;
        RECT 1.250 0.480 1.555 1.010 ;
        RECT 2.165 0.480 2.415 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.105 2.440 0.435 2.980 ;
        RECT 0.620 2.610 0.950 3.245 ;
        RECT 1.520 2.610 1.850 3.245 ;
        RECT 2.420 2.610 2.750 3.245 ;
        RECT 2.940 2.905 4.090 3.075 ;
        RECT 0.105 2.270 2.640 2.440 ;
        RECT 0.105 1.275 0.435 2.270 ;
        RECT 2.470 2.020 2.640 2.270 ;
        RECT 2.940 2.190 3.270 2.905 ;
        RECT 2.470 1.850 3.290 2.020 ;
        RECT 1.590 1.350 2.755 1.680 ;
        RECT 2.960 1.450 3.290 1.850 ;
        RECT 2.585 1.280 2.755 1.350 ;
        RECT 3.470 1.280 3.720 2.735 ;
        RECT 3.920 2.120 4.090 2.905 ;
        RECT 4.290 2.290 4.540 3.245 ;
        RECT 4.740 2.120 5.070 2.980 ;
        RECT 5.270 2.290 5.520 3.245 ;
        RECT 5.720 2.120 5.970 2.980 ;
        RECT 3.920 1.950 5.970 2.120 ;
        RECT 3.920 1.940 4.090 1.950 ;
        RECT 5.720 1.940 5.970 1.950 ;
        RECT 0.105 0.840 0.615 1.275 ;
        RECT 0.795 0.085 1.045 1.275 ;
        RECT 2.585 1.110 5.035 1.280 ;
        RECT 1.735 0.085 1.985 0.840 ;
        RECT 2.595 0.085 2.845 0.940 ;
        RECT 3.085 0.595 3.415 1.110 ;
        RECT 3.595 0.085 3.765 0.940 ;
        RECT 4.435 0.425 4.605 0.940 ;
        RECT 4.785 0.595 5.035 1.110 ;
        RECT 5.215 0.425 5.545 1.275 ;
        RECT 4.435 0.255 5.545 0.425 ;
        RECT 5.725 0.085 5.975 1.275 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__a21bo_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a21boi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21boi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.295 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.180 3.235 1.550 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.255 0.450 1.605 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.530 0.245 3.070 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.515200 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.920 1.525 2.980 ;
        RECT 1.275 1.890 1.525 1.920 ;
        RECT 1.275 1.720 1.875 1.890 ;
        RECT 1.705 1.180 1.875 1.720 ;
        RECT 1.705 1.010 2.060 1.180 ;
        RECT 1.810 0.350 2.060 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.105 1.945 0.435 2.980 ;
        RECT 0.635 2.115 0.885 3.245 ;
        RECT 1.725 2.230 2.020 2.980 ;
        RECT 2.190 2.400 2.520 3.245 ;
        RECT 2.690 2.230 2.985 2.980 ;
        RECT 1.725 2.060 2.985 2.230 ;
        RECT 0.105 1.775 0.915 1.945 ;
        RECT 2.655 1.820 2.985 2.060 ;
        RECT 0.745 1.550 0.915 1.775 ;
        RECT 0.745 1.220 1.535 1.550 ;
        RECT 0.745 1.050 0.950 1.220 ;
        RECT 0.620 0.540 0.950 1.050 ;
        RECT 1.120 0.760 1.450 1.050 ;
        RECT 1.120 0.085 1.630 0.760 ;
        RECT 2.630 0.085 2.960 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a21boi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21boi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.320 2.815 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.265 1.220 3.715 1.550 ;
        RECT 3.485 1.180 3.715 1.220 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.475 1.780 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.180 0.245 4.280 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.750400 ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.410 1.945 2.735 ;
        RECT 1.615 1.150 2.275 1.410 ;
        RECT 1.270 0.980 2.900 1.150 ;
        RECT 1.270 0.350 1.440 0.980 ;
        RECT 2.570 0.770 2.900 0.980 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.195 1.950 0.445 3.245 ;
        RECT 0.645 1.940 0.975 2.980 ;
        RECT 0.805 1.650 0.975 1.940 ;
        RECT 1.165 2.905 2.315 3.075 ;
        RECT 1.165 1.820 1.415 2.905 ;
        RECT 2.115 2.120 2.315 2.905 ;
        RECT 2.515 2.290 2.845 3.245 ;
        RECT 3.045 2.120 3.215 2.980 ;
        RECT 2.115 1.950 3.215 2.120 ;
        RECT 3.415 2.060 3.765 3.245 ;
        RECT 2.115 1.820 2.315 1.950 ;
        RECT 3.045 1.890 3.215 1.950 ;
        RECT 3.965 1.890 4.215 2.980 ;
        RECT 3.045 1.720 4.215 1.890 ;
        RECT 0.805 1.320 1.395 1.650 ;
        RECT 0.805 1.280 0.975 1.320 ;
        RECT 0.270 1.110 0.975 1.280 ;
        RECT 0.270 0.450 0.520 1.110 ;
        RECT 3.080 1.010 3.250 1.050 ;
        RECT 3.940 1.010 4.190 1.130 ;
        RECT 0.760 0.085 1.090 0.940 ;
        RECT 3.080 0.840 4.190 1.010 ;
        RECT 1.620 0.085 1.950 0.810 ;
        RECT 3.080 0.600 3.250 0.840 ;
        RECT 2.140 0.350 3.250 0.600 ;
        RECT 3.430 0.085 3.760 0.670 ;
        RECT 3.940 0.350 4.190 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a21boi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21boi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.430 1.795 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.430 3.715 1.780 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.490 7.555 1.820 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.245 6.750 1.240 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.500800 ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.990 4.495 2.735 ;
        RECT 5.065 1.990 5.395 2.735 ;
        RECT 4.165 1.820 5.395 1.990 ;
        RECT 4.165 1.780 4.745 1.820 ;
        RECT 3.965 1.260 4.745 1.780 ;
        RECT 1.480 1.150 4.745 1.260 ;
        RECT 0.700 0.940 0.950 1.130 ;
        RECT 1.480 1.090 5.720 1.150 ;
        RECT 1.480 0.940 1.810 1.090 ;
        RECT 4.575 0.980 5.720 1.090 ;
        RECT 0.700 0.770 1.810 0.940 ;
        RECT 4.610 0.350 4.860 0.980 ;
        RECT 5.470 0.350 5.720 0.980 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.115 2.120 0.365 2.980 ;
        RECT 0.565 2.290 0.895 3.245 ;
        RECT 1.095 2.120 1.265 2.980 ;
        RECT 1.465 2.290 1.795 3.245 ;
        RECT 1.995 2.120 2.165 2.980 ;
        RECT 2.365 2.290 2.615 3.245 ;
        RECT 2.815 2.120 3.145 2.980 ;
        RECT 3.345 2.290 3.515 3.245 ;
        RECT 3.715 2.905 5.845 3.075 ;
        RECT 3.715 2.120 3.995 2.905 ;
        RECT 4.665 2.160 4.895 2.905 ;
        RECT 0.115 1.950 3.995 2.120 ;
        RECT 1.995 1.820 2.165 1.950 ;
        RECT 5.565 1.820 5.845 2.905 ;
        RECT 6.035 2.330 6.365 3.245 ;
        RECT 6.535 2.160 6.815 2.980 ;
        RECT 6.025 1.990 6.815 2.160 ;
        RECT 7.015 2.100 7.265 3.245 ;
        RECT 6.025 1.650 6.195 1.990 ;
        RECT 4.915 1.320 6.195 1.650 ;
        RECT 6.025 1.150 6.660 1.320 ;
        RECT 0.190 0.600 0.520 1.130 ;
        RECT 1.990 0.750 3.960 0.920 ;
        RECT 1.990 0.600 2.160 0.750 ;
        RECT 0.190 0.350 2.160 0.600 ;
        RECT 2.340 0.085 2.670 0.580 ;
        RECT 2.850 0.510 3.020 0.750 ;
        RECT 3.200 0.085 3.530 0.580 ;
        RECT 3.710 0.510 3.960 0.750 ;
        RECT 4.180 0.085 4.430 0.880 ;
        RECT 5.040 0.085 5.290 0.810 ;
        RECT 5.900 0.085 6.230 0.980 ;
        RECT 6.400 0.350 6.660 1.150 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__a21boi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.450 2.375 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 0.570 3.235 0.670 ;
        RECT 2.645 0.255 3.235 0.570 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.450 1.835 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.735 0.245 3.130 1.450 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.435 2.980 ;
        RECT 0.085 1.150 0.255 1.820 ;
        RECT 0.085 0.980 1.075 1.150 ;
        RECT 0.825 0.670 1.075 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.635 1.820 0.885 3.245 ;
        RECT 1.245 1.950 1.605 2.980 ;
        RECT 1.805 2.120 2.135 2.980 ;
        RECT 2.335 2.290 2.535 3.245 ;
        RECT 2.735 2.120 3.065 2.980 ;
        RECT 1.805 1.950 3.065 2.120 ;
        RECT 1.245 1.650 1.415 1.950 ;
        RECT 2.735 1.940 3.065 1.950 ;
        RECT 0.425 1.320 1.415 1.650 ;
        RECT 1.245 1.280 1.415 1.320 ;
        RECT 1.245 1.110 2.135 1.280 ;
        RECT 1.255 0.085 1.585 0.940 ;
        RECT 1.805 0.660 2.135 1.110 ;
        RECT 2.710 1.010 3.040 1.340 ;
        RECT 2.305 0.840 3.040 1.010 ;
        RECT 2.305 0.085 2.475 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a21o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.200 1.180 2.755 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.180 3.255 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.180 1.990 1.535 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.205 0.245 3.305 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.570 1.890 0.850 2.980 ;
        RECT 0.570 1.550 0.900 1.890 ;
        RECT 0.725 1.050 0.900 1.550 ;
        RECT 0.725 0.350 1.055 1.050 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.120 1.820 0.370 3.245 ;
        RECT 1.020 2.045 1.350 3.245 ;
        RECT 1.540 1.875 1.790 2.980 ;
        RECT 1.070 1.705 1.790 1.875 ;
        RECT 1.990 1.890 2.240 2.980 ;
        RECT 2.440 2.060 2.770 3.245 ;
        RECT 2.970 1.890 3.220 2.980 ;
        RECT 1.990 1.720 3.220 1.890 ;
        RECT 1.070 1.220 1.395 1.705 ;
        RECT 0.295 0.085 0.545 1.130 ;
        RECT 1.225 1.010 1.395 1.220 ;
        RECT 1.225 0.840 2.295 1.010 ;
        RECT 1.225 0.085 1.795 0.670 ;
        RECT 1.965 0.350 2.295 0.840 ;
        RECT 2.865 0.085 3.195 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a21o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.450 4.195 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.260 4.905 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.425 1.435 2.755 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 1.140 3.210 1.240 ;
        RECT 0.040 0.245 5.600 1.140 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.685 1.970 0.855 2.980 ;
        RECT 1.505 1.970 1.835 2.980 ;
        RECT 0.125 1.800 1.835 1.970 ;
        RECT 0.125 1.130 0.355 1.800 ;
        RECT 0.125 0.960 1.690 1.130 ;
        RECT 0.660 0.350 0.830 0.960 ;
        RECT 1.440 0.350 1.690 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.155 2.140 0.485 3.245 ;
        RECT 1.055 2.140 1.305 3.245 ;
        RECT 2.035 1.950 2.285 3.245 ;
        RECT 2.475 2.905 3.625 3.075 ;
        RECT 2.475 1.950 2.725 2.905 ;
        RECT 0.635 1.300 2.205 1.630 ;
        RECT 1.870 1.265 2.205 1.300 ;
        RECT 2.925 1.280 3.255 2.735 ;
        RECT 3.455 2.120 3.625 2.905 ;
        RECT 3.825 2.290 4.075 3.245 ;
        RECT 4.275 2.120 4.525 2.980 ;
        RECT 4.725 2.290 5.055 3.245 ;
        RECT 5.255 2.120 5.505 2.980 ;
        RECT 3.455 1.950 5.505 2.120 ;
        RECT 5.255 1.940 5.505 1.950 ;
        RECT 2.925 1.265 4.220 1.280 ;
        RECT 1.870 1.110 4.220 1.265 ;
        RECT 1.870 1.095 3.255 1.110 ;
        RECT 0.150 0.085 0.480 0.790 ;
        RECT 1.010 0.085 1.260 0.790 ;
        RECT 1.870 0.085 2.120 0.925 ;
        RECT 2.360 0.450 2.610 1.095 ;
        RECT 2.790 0.085 3.120 0.925 ;
        RECT 3.460 0.425 3.790 0.940 ;
        RECT 3.960 0.595 4.220 1.110 ;
        RECT 4.400 0.920 5.510 1.090 ;
        RECT 4.400 0.425 4.570 0.920 ;
        RECT 3.460 0.255 4.570 0.425 ;
        RECT 4.750 0.085 5.080 0.750 ;
        RECT 5.260 0.350 5.510 0.920 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__a21o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 1.050 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.560 1.190 1.815 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.245 1.900 1.240 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596600 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.890 1.815 2.980 ;
        RECT 1.220 1.720 1.815 1.890 ;
        RECT 1.220 1.180 1.390 1.720 ;
        RECT 0.920 1.010 1.390 1.180 ;
        RECT 0.920 0.350 1.290 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.105 2.230 0.400 2.980 ;
        RECT 0.570 2.400 0.900 3.245 ;
        RECT 1.070 2.230 1.365 2.980 ;
        RECT 0.105 2.060 1.365 2.230 ;
        RECT 0.105 1.985 0.955 2.060 ;
        RECT 0.105 1.820 0.435 1.985 ;
        RECT 0.130 0.085 0.460 1.010 ;
        RECT 1.560 0.085 1.790 1.020 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__a21oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 3.350 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.755 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.435 0.435 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.270 1.405 1.780 1.450 ;
        RECT 1.270 1.240 2.255 1.405 ;
        RECT 0.010 0.245 3.780 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.739300 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.780 1.395 2.735 ;
        RECT 0.605 1.550 1.395 1.780 ;
        RECT 0.605 0.920 0.860 1.550 ;
        RECT 2.930 0.920 3.180 1.130 ;
        RECT 0.605 0.750 3.180 0.920 ;
        RECT 0.605 0.350 0.860 0.750 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.615 2.905 1.845 3.075 ;
        RECT 0.615 1.950 0.895 2.905 ;
        RECT 1.565 2.460 1.845 2.905 ;
        RECT 2.045 2.630 2.305 3.245 ;
        RECT 2.475 2.460 2.805 2.980 ;
        RECT 3.005 2.630 3.175 3.245 ;
        RECT 3.375 2.460 3.705 2.980 ;
        RECT 1.565 2.290 3.705 2.460 ;
        RECT 1.565 1.950 3.690 2.120 ;
        RECT 1.565 1.260 1.775 1.950 ;
        RECT 0.100 0.085 0.430 1.130 ;
        RECT 1.360 1.090 1.775 1.260 ;
        RECT 3.520 1.130 3.690 1.950 ;
        RECT 3.360 0.580 3.690 1.130 ;
        RECT 2.000 0.085 2.330 0.580 ;
        RECT 2.500 0.330 3.690 0.580 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a21oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a21oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.350 3.935 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.785 1.350 2.275 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 4.235 1.350 5.245 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.290 0.245 5.680 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.478600 ;
    PORT
      LAYER li1 ;
        RECT 4.355 2.120 4.685 2.735 ;
        RECT 5.255 2.120 5.585 2.735 ;
        RECT 2.525 1.950 5.585 2.120 ;
        RECT 2.525 1.180 2.755 1.950 ;
        RECT 2.525 1.010 5.590 1.180 ;
        RECT 2.525 0.880 4.650 1.010 ;
        RECT 2.525 0.595 2.780 0.880 ;
        RECT 4.400 0.350 4.650 0.880 ;
        RECT 5.340 0.350 5.590 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.305 2.120 0.555 2.980 ;
        RECT 0.755 2.290 1.005 3.245 ;
        RECT 1.205 2.120 1.535 2.980 ;
        RECT 1.735 2.290 1.905 3.245 ;
        RECT 2.105 2.460 2.355 2.980 ;
        RECT 2.555 2.630 2.805 3.245 ;
        RECT 3.005 2.460 3.335 2.980 ;
        RECT 3.535 2.630 3.705 3.245 ;
        RECT 3.905 2.905 6.035 3.075 ;
        RECT 3.905 2.460 4.155 2.905 ;
        RECT 2.105 2.290 4.155 2.460 ;
        RECT 4.885 2.290 5.055 2.905 ;
        RECT 2.105 2.120 2.355 2.290 ;
        RECT 0.305 1.950 2.355 2.120 ;
        RECT 0.305 1.820 0.555 1.950 ;
        RECT 5.785 1.820 6.035 2.905 ;
        RECT 0.380 1.010 2.350 1.180 ;
        RECT 0.380 0.350 0.630 1.010 ;
        RECT 0.810 0.085 1.140 0.840 ;
        RECT 1.320 0.350 1.490 1.010 ;
        RECT 1.670 0.085 2.000 0.840 ;
        RECT 2.180 0.425 2.350 1.010 ;
        RECT 2.960 0.425 3.290 0.710 ;
        RECT 3.820 0.425 4.150 0.710 ;
        RECT 2.180 0.255 4.150 0.425 ;
        RECT 4.830 0.085 5.160 0.840 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__a21oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a22o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.350 2.295 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.505 0.355 0.670 ;
        RECT 0.125 0.255 0.560 0.505 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.425 1.470 1.795 1.800 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.470 1.215 1.800 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130 1.165 1.055 1.385 ;
        RECT 2.405 1.165 3.345 1.240 ;
        RECT 0.130 0.245 3.345 1.165 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 2.925 0.350 3.255 2.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.195 1.970 0.445 3.245 ;
        RECT 0.645 2.905 1.995 3.075 ;
        RECT 0.645 1.970 0.895 2.905 ;
        RECT 1.095 2.140 1.425 2.735 ;
        RECT 1.595 2.310 1.995 2.905 ;
        RECT 2.165 2.310 2.725 3.245 ;
        RECT 1.095 1.970 2.755 2.140 ;
        RECT 0.220 1.130 1.285 1.300 ;
        RECT 2.505 1.180 2.755 1.970 ;
        RECT 0.220 0.840 0.550 1.130 ;
        RECT 0.730 0.085 0.945 0.960 ;
        RECT 1.115 0.625 1.285 1.130 ;
        RECT 1.485 1.010 2.755 1.180 ;
        RECT 1.485 0.795 1.815 1.010 ;
        RECT 1.115 0.375 2.245 0.625 ;
        RECT 2.495 0.085 2.745 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a22o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a22o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a22o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.350 1.905 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.350 3.735 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.350 2.495 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.705 1.350 3.235 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 3.810 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.905 2.290 1.185 2.980 ;
        RECT 0.905 1.890 1.075 2.290 ;
        RECT 0.530 1.720 1.075 1.890 ;
        RECT 0.530 0.350 0.860 1.720 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.485 2.060 0.735 3.245 ;
        RECT 1.385 2.290 1.715 3.245 ;
        RECT 1.925 2.905 3.225 3.075 ;
        RECT 1.925 2.290 2.255 2.905 ;
        RECT 2.455 2.120 2.705 2.735 ;
        RECT 1.245 1.950 2.705 2.120 ;
        RECT 2.875 1.950 3.225 2.905 ;
        RECT 3.395 1.950 3.725 3.245 ;
        RECT 1.245 1.550 1.415 1.950 ;
        RECT 1.085 1.180 1.415 1.550 ;
        RECT 0.100 0.085 0.350 1.130 ;
        RECT 1.085 1.010 2.330 1.180 ;
        RECT 1.040 0.085 1.290 0.840 ;
        RECT 1.500 0.425 1.830 0.840 ;
        RECT 2.000 0.595 2.330 1.010 ;
        RECT 2.500 1.010 3.700 1.180 ;
        RECT 2.500 0.425 2.670 1.010 ;
        RECT 1.500 0.255 2.670 0.425 ;
        RECT 2.870 0.085 3.200 0.840 ;
        RECT 3.370 0.350 3.700 1.010 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a22o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a22o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.450 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.955 0.505 5.125 0.670 ;
        RECT 4.955 0.255 5.320 0.505 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.495 1.435 3.825 1.765 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.935 4.195 2.150 ;
        RECT 3.155 1.765 3.325 1.935 ;
        RECT 3.025 1.435 3.325 1.765 ;
        RECT 4.025 1.770 4.195 1.935 ;
        RECT 4.025 1.440 4.655 1.770 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.030 1.370 7.005 1.385 ;
        RECT 0.885 0.245 7.005 1.370 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.705 1.650 0.875 2.980 ;
        RECT 1.525 1.650 1.855 2.980 ;
        RECT 0.705 1.410 1.855 1.650 ;
        RECT 0.125 1.180 1.855 1.410 ;
        RECT 0.125 1.140 2.515 1.180 ;
        RECT 1.405 1.010 2.515 1.140 ;
        RECT 1.405 0.480 1.655 1.010 ;
        RECT 2.265 0.480 2.515 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.175 1.900 0.505 3.245 ;
        RECT 1.075 1.820 1.325 3.245 ;
        RECT 2.055 1.850 2.305 3.245 ;
        RECT 2.475 2.980 3.515 3.075 ;
        RECT 2.475 2.905 4.415 2.980 ;
        RECT 2.475 1.680 2.645 2.905 ;
        RECT 2.815 2.490 2.985 2.735 ;
        RECT 3.185 2.660 4.415 2.905 ;
        RECT 4.615 2.490 4.865 2.980 ;
        RECT 2.815 2.320 4.865 2.490 ;
        RECT 2.815 1.940 2.985 2.320 ;
        RECT 4.615 2.120 4.865 2.320 ;
        RECT 5.035 2.290 5.510 3.245 ;
        RECT 5.680 2.120 5.930 2.980 ;
        RECT 6.130 2.290 6.460 3.245 ;
        RECT 6.660 2.120 6.910 2.980 ;
        RECT 4.615 1.950 6.910 2.120 ;
        RECT 4.615 1.940 4.865 1.950 ;
        RECT 6.660 1.940 6.910 1.950 ;
        RECT 2.025 1.350 2.855 1.680 ;
        RECT 2.685 1.265 2.855 1.350 ;
        RECT 5.725 1.265 6.055 1.275 ;
        RECT 2.685 1.095 6.055 1.265 ;
        RECT 3.630 1.000 3.960 1.095 ;
        RECT 5.725 1.015 6.055 1.095 ;
        RECT 0.975 0.085 1.225 0.970 ;
        RECT 1.835 0.085 2.085 0.840 ;
        RECT 2.695 0.085 3.025 0.925 ;
        RECT 4.140 0.830 4.355 0.925 ;
        RECT 3.200 0.580 4.355 0.830 ;
        RECT 4.535 0.085 4.785 0.925 ;
        RECT 6.235 0.845 6.405 1.275 ;
        RECT 5.295 0.675 6.405 0.845 ;
        RECT 6.235 0.595 6.405 0.675 ;
        RECT 6.585 0.085 6.915 1.275 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__a22o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a22oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.755 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.350 1.335 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.250 0.245 2.630 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.624600 ;
    PORT
      LAYER li1 ;
        RECT 0.845 2.120 1.015 2.735 ;
        RECT 0.605 1.950 1.015 2.120 ;
        RECT 0.605 1.180 0.835 1.950 ;
        RECT 0.605 1.010 1.570 1.180 ;
        RECT 1.130 0.350 1.570 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.315 2.905 1.545 3.075 ;
        RECT 0.315 2.290 0.645 2.905 ;
        RECT 1.215 2.120 1.545 2.905 ;
        RECT 1.715 2.290 2.065 3.245 ;
        RECT 2.235 2.120 2.565 2.980 ;
        RECT 1.215 1.950 2.565 2.120 ;
        RECT 0.340 0.085 0.670 0.840 ;
        RECT 2.210 0.085 2.540 1.130 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__a22oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a22oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.710 1.950 2.210 2.120 ;
        RECT 0.710 1.780 0.880 1.950 ;
        RECT 0.125 1.430 0.880 1.780 ;
        RECT 1.880 1.430 2.210 1.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.430 1.420 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.720 1.260 3.235 1.550 ;
        RECT 3.905 1.300 4.370 1.630 ;
        RECT 3.905 1.260 4.075 1.300 ;
        RECT 2.720 1.090 4.075 1.260 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.430 3.735 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.195 0.245 4.585 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.497400 ;
    PORT
      LAYER li1 ;
        RECT 2.930 2.120 3.130 2.735 ;
        RECT 3.860 2.120 4.030 2.735 ;
        RECT 2.930 1.950 4.710 2.120 ;
        RECT 2.930 1.890 3.130 1.950 ;
        RECT 2.380 1.720 3.130 1.890 ;
        RECT 2.380 1.260 2.550 1.720 ;
        RECT 0.285 1.090 2.550 1.260 ;
        RECT 4.540 1.130 4.710 1.950 ;
        RECT 0.285 0.350 0.535 1.090 ;
        RECT 2.040 0.810 2.550 1.090 ;
        RECT 2.145 0.350 2.550 0.810 ;
        RECT 4.245 0.350 4.710 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.290 2.460 0.540 2.980 ;
        RECT 0.740 2.630 0.990 3.245 ;
        RECT 1.190 2.460 1.520 2.980 ;
        RECT 1.690 2.630 2.230 3.245 ;
        RECT 2.400 2.905 4.560 3.075 ;
        RECT 2.400 2.460 2.730 2.905 ;
        RECT 0.290 2.290 2.730 2.460 ;
        RECT 3.330 2.290 3.660 2.905 ;
        RECT 4.230 2.290 4.560 2.905 ;
        RECT 0.290 1.950 0.540 2.290 ;
        RECT 2.400 2.060 2.730 2.290 ;
        RECT 0.715 0.750 1.815 0.920 ;
        RECT 0.715 0.330 0.965 0.750 ;
        RECT 1.645 0.640 1.815 0.750 ;
        RECT 2.835 0.750 4.065 0.920 ;
        RECT 1.145 0.085 1.475 0.580 ;
        RECT 1.645 0.350 1.975 0.640 ;
        RECT 2.835 0.330 3.135 0.750 ;
        RECT 3.305 0.085 3.635 0.580 ;
        RECT 3.815 0.330 4.065 0.750 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__a22oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a22oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 5.635 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.350 7.465 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.350 3.275 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 1.955 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.110 0.245 8.020 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.172800 ;
    PORT
      LAYER li1 ;
        RECT 0.635 2.120 0.885 2.735 ;
        RECT 1.615 2.120 1.785 2.735 ;
        RECT 2.515 2.120 2.685 2.735 ;
        RECT 3.415 2.120 3.615 2.735 ;
        RECT 0.635 1.950 3.615 2.120 ;
        RECT 3.445 1.520 3.615 1.950 ;
        RECT 3.445 1.180 4.195 1.520 ;
        RECT 2.350 1.130 4.195 1.180 ;
        RECT 2.350 1.010 5.780 1.130 ;
        RECT 2.350 0.595 2.680 1.010 ;
        RECT 3.210 0.850 5.780 1.010 ;
        RECT 3.210 0.770 3.990 0.850 ;
        RECT 5.450 0.770 5.780 0.850 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.185 2.905 4.035 3.075 ;
        RECT 0.185 1.820 0.435 2.905 ;
        RECT 1.085 2.290 1.415 2.905 ;
        RECT 1.985 2.290 2.315 2.905 ;
        RECT 2.885 2.290 3.215 2.905 ;
        RECT 3.785 2.120 4.035 2.905 ;
        RECT 4.235 2.290 4.565 3.245 ;
        RECT 4.765 2.120 5.015 2.980 ;
        RECT 5.185 2.290 5.645 3.245 ;
        RECT 5.815 2.120 6.065 2.980 ;
        RECT 6.265 2.290 6.595 3.245 ;
        RECT 6.795 2.120 6.965 2.980 ;
        RECT 7.165 2.290 7.495 3.245 ;
        RECT 7.695 2.120 7.945 2.980 ;
        RECT 3.785 1.950 7.945 2.120 ;
        RECT 3.785 1.820 4.035 1.950 ;
        RECT 7.695 1.820 7.945 1.950 ;
        RECT 0.200 1.010 2.170 1.180 ;
        RECT 0.200 0.350 0.450 1.010 ;
        RECT 0.630 0.085 0.880 0.840 ;
        RECT 1.060 0.350 1.310 1.010 ;
        RECT 1.490 0.085 1.820 0.840 ;
        RECT 2.000 0.425 2.170 1.010 ;
        RECT 5.960 1.010 7.930 1.180 ;
        RECT 2.860 0.600 3.030 0.840 ;
        RECT 4.160 0.600 4.490 0.680 ;
        RECT 5.960 0.600 6.130 1.010 ;
        RECT 2.860 0.425 3.970 0.600 ;
        RECT 2.000 0.255 3.970 0.425 ;
        RECT 4.160 0.350 6.130 0.600 ;
        RECT 6.310 0.085 6.560 0.840 ;
        RECT 6.740 0.350 6.990 1.010 ;
        RECT 7.170 0.085 7.420 0.840 ;
        RECT 7.600 0.350 7.930 1.010 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__a22oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.490 2.405 1.800 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.490 1.865 1.800 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.490 1.325 1.800 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.255 2.815 0.640 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.695 1.370 3.210 1.385 ;
        RECT 0.040 0.245 3.210 1.370 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.850 0.435 2.980 ;
        RECT 0.085 1.180 0.255 1.850 ;
        RECT 0.085 0.480 0.450 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.605 1.970 1.065 3.245 ;
        RECT 1.235 2.140 1.565 2.980 ;
        RECT 1.735 2.310 2.145 3.245 ;
        RECT 2.315 2.140 2.645 2.980 ;
        RECT 1.235 1.970 2.645 2.140 ;
        RECT 0.425 1.350 0.825 1.680 ;
        RECT 0.620 1.320 0.825 1.350 ;
        RECT 2.845 1.320 3.095 2.980 ;
        RECT 0.620 1.150 3.095 1.320 ;
        RECT 0.620 0.085 1.200 0.980 ;
        RECT 2.280 0.810 2.610 1.150 ;
        RECT 2.790 0.810 3.155 0.980 ;
        RECT 2.985 0.085 3.155 0.810 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a31o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a31o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.665 1.180 3.235 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.425 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.180 1.855 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.180 3.735 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.800 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.820 0.920 2.980 ;
        RECT 0.615 1.130 0.785 1.820 ;
        RECT 0.615 0.350 0.890 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.185 1.820 0.435 3.245 ;
        RECT 1.090 2.060 1.625 3.245 ;
        RECT 1.795 2.230 2.125 2.860 ;
        RECT 2.350 2.400 2.680 3.245 ;
        RECT 2.885 2.230 3.215 2.860 ;
        RECT 1.795 2.060 3.215 2.230 ;
        RECT 3.385 1.890 3.725 2.860 ;
        RECT 1.135 1.720 3.725 1.890 ;
        RECT 1.135 1.630 1.305 1.720 ;
        RECT 0.955 1.300 1.305 1.630 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 1.135 1.010 1.305 1.300 ;
        RECT 1.135 0.840 3.180 1.010 ;
        RECT 1.060 0.085 1.730 0.600 ;
        RECT 2.850 0.350 3.180 0.840 ;
        RECT 3.360 0.085 3.690 1.010 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a31o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.450 4.675 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.450 5.865 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.115 1.450 7.075 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.565 1.470 3.235 1.800 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 2.370 1.240 ;
        RECT 0.005 0.245 7.140 1.140 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.138200 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.890 0.895 2.980 ;
        RECT 1.565 1.890 1.895 2.980 ;
        RECT 0.565 1.720 1.895 1.890 ;
        RECT 0.565 1.550 0.895 1.720 ;
        RECT 0.615 1.000 0.865 1.550 ;
        RECT 0.615 0.830 1.725 1.000 ;
        RECT 0.615 0.350 0.865 0.830 ;
        RECT 1.555 0.330 1.725 0.830 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.065 2.060 1.395 3.245 ;
        RECT 2.065 1.820 2.395 3.245 ;
        RECT 2.625 2.810 4.075 2.980 ;
        RECT 2.625 1.970 2.955 2.810 ;
        RECT 3.125 1.970 3.575 2.640 ;
        RECT 1.065 1.300 2.335 1.550 ;
        RECT 3.405 1.300 3.575 1.970 ;
        RECT 3.745 2.120 4.075 2.810 ;
        RECT 4.245 2.290 4.575 3.245 ;
        RECT 4.745 2.120 5.075 2.980 ;
        RECT 5.245 2.290 5.575 3.245 ;
        RECT 5.755 2.120 6.085 2.980 ;
        RECT 6.255 2.290 6.585 3.245 ;
        RECT 6.755 2.120 7.085 2.980 ;
        RECT 3.745 1.950 7.085 2.120 ;
        RECT 1.065 1.280 3.590 1.300 ;
        RECT 1.065 1.220 4.750 1.280 ;
        RECT 1.895 1.130 4.750 1.220 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 1.045 0.085 1.375 0.660 ;
        RECT 1.930 0.085 2.260 0.960 ;
        RECT 2.490 0.350 2.740 1.130 ;
        RECT 3.420 1.110 4.750 1.130 ;
        RECT 2.920 0.085 3.250 0.960 ;
        RECT 3.420 0.350 3.750 1.110 ;
        RECT 3.920 0.425 4.250 0.940 ;
        RECT 4.420 0.595 4.750 1.110 ;
        RECT 4.980 1.110 7.030 1.280 ;
        RECT 4.980 0.595 5.230 1.110 ;
        RECT 5.410 0.425 5.740 0.940 ;
        RECT 3.920 0.255 5.740 0.425 ;
        RECT 5.920 0.350 6.090 1.110 ;
        RECT 6.270 0.085 6.600 0.940 ;
        RECT 6.780 0.350 7.030 1.110 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__a31o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a31oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.180 1.865 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.810 1.315 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.455 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.775 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.245 2.670 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641200 ;
    PORT
      LAYER li1 ;
        RECT 2.255 1.890 2.755 2.980 ;
        RECT 0.625 1.720 2.755 1.890 ;
        RECT 0.625 0.520 0.795 1.720 ;
        RECT 1.730 0.520 2.060 1.010 ;
        RECT 0.625 0.350 2.060 0.520 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.125 1.820 0.455 3.245 ;
        RECT 0.665 2.230 0.995 2.980 ;
        RECT 1.205 2.400 1.535 3.245 ;
        RECT 1.755 2.230 2.085 2.980 ;
        RECT 0.665 2.060 2.085 2.230 ;
        RECT 0.125 0.085 0.455 1.010 ;
        RECT 2.230 0.085 2.560 1.010 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__a31oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.505 1.430 4.195 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.430 1.545 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.260 0.435 1.550 ;
        RECT 1.785 1.260 2.115 1.550 ;
        RECT 0.105 1.090 2.115 1.260 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.180 2.995 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.090800 ;
    PORT
      LAYER li1 ;
        RECT 2.475 1.890 2.805 2.735 ;
        RECT 2.475 1.720 3.335 1.890 ;
        RECT 3.165 1.260 3.335 1.720 ;
        RECT 3.165 1.090 4.205 1.260 ;
        RECT 2.545 0.425 3.260 0.580 ;
        RECT 3.875 0.425 4.205 1.090 ;
        RECT 2.545 0.255 4.205 0.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.120 0.365 2.980 ;
        RECT 0.565 2.290 0.895 3.245 ;
        RECT 1.065 2.120 1.395 2.980 ;
        RECT 1.595 2.290 1.845 3.245 ;
        RECT 2.015 2.905 3.255 3.075 ;
        RECT 2.015 2.120 2.275 2.905 ;
        RECT 0.115 1.950 2.275 2.120 ;
        RECT 2.975 2.230 3.255 2.905 ;
        RECT 3.425 2.400 3.755 3.245 ;
        RECT 3.925 2.230 4.205 2.980 ;
        RECT 2.975 2.060 4.205 2.230 ;
        RECT 3.875 1.950 4.205 2.060 ;
        RECT 0.115 1.820 0.365 1.950 ;
        RECT 0.115 0.085 0.365 0.920 ;
        RECT 0.545 0.425 0.875 0.920 ;
        RECT 1.045 0.750 3.705 0.920 ;
        RECT 1.045 0.595 1.375 0.750 ;
        RECT 3.430 0.670 3.705 0.750 ;
        RECT 1.545 0.425 1.875 0.580 ;
        RECT 0.545 0.255 1.875 0.425 ;
        RECT 2.045 0.085 2.375 0.580 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a31oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.350 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.350 4.195 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.745 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.350 8.515 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 8.635 1.240 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.621350 ;
    PORT
      LAYER li1 ;
        RECT 6.845 2.120 7.175 2.735 ;
        RECT 7.745 2.120 8.075 2.735 ;
        RECT 4.445 1.950 8.075 2.120 ;
        RECT 4.445 1.180 4.690 1.950 ;
        RECT 4.445 1.130 8.525 1.180 ;
        RECT 4.350 1.010 8.525 1.130 ;
        RECT 4.350 0.965 5.840 1.010 ;
        RECT 4.350 0.770 4.685 0.965 ;
        RECT 5.510 0.595 5.840 0.965 ;
        RECT 6.510 0.350 6.840 1.010 ;
        RECT 8.195 0.350 8.525 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.115 2.120 0.395 2.980 ;
        RECT 0.565 2.290 0.895 3.245 ;
        RECT 1.065 2.120 1.295 2.935 ;
        RECT 1.465 2.290 1.795 3.245 ;
        RECT 1.965 2.150 2.195 2.950 ;
        RECT 2.365 2.320 2.695 3.245 ;
        RECT 2.865 2.150 3.195 2.980 ;
        RECT 3.365 2.290 3.695 3.245 ;
        RECT 3.865 2.460 4.195 2.980 ;
        RECT 4.365 2.630 4.695 3.245 ;
        RECT 4.865 2.460 5.675 2.930 ;
        RECT 5.845 2.630 6.175 3.245 ;
        RECT 6.345 2.905 8.525 3.075 ;
        RECT 6.345 2.460 6.675 2.905 ;
        RECT 3.865 2.290 6.675 2.460 ;
        RECT 7.375 2.290 7.575 2.905 ;
        RECT 1.965 2.120 3.195 2.150 ;
        RECT 3.865 2.120 4.195 2.290 ;
        RECT 0.115 1.950 4.195 2.120 ;
        RECT 8.255 1.950 8.525 2.905 ;
        RECT 1.915 1.820 2.245 1.950 ;
        RECT 0.130 1.010 4.120 1.180 ;
        RECT 0.130 0.350 0.380 1.010 ;
        RECT 0.560 0.085 0.890 0.840 ;
        RECT 1.070 0.350 1.240 1.010 ;
        RECT 1.420 0.085 1.750 0.840 ;
        RECT 1.920 0.330 2.170 1.010 ;
        RECT 2.350 0.425 2.655 0.840 ;
        RECT 2.825 0.595 3.120 1.010 ;
        RECT 3.290 0.425 3.620 0.840 ;
        RECT 3.790 0.595 4.120 1.010 ;
        RECT 4.935 0.425 5.265 0.795 ;
        RECT 6.010 0.425 6.340 0.840 ;
        RECT 2.350 0.255 6.340 0.425 ;
        RECT 7.010 0.085 8.025 0.840 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__a31oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a32o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a32o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.190 2.375 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.190 1.835 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.190 1.315 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.190 3.005 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.290 1.210 3.715 1.550 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.810 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.455 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.445 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.625 2.060 1.015 3.245 ;
        RECT 1.205 2.230 1.535 2.860 ;
        RECT 1.800 2.400 2.130 3.245 ;
        RECT 2.395 2.905 3.725 3.075 ;
        RECT 2.395 2.230 2.725 2.905 ;
        RECT 1.205 2.060 2.725 2.230 ;
        RECT 2.895 1.890 3.225 2.735 ;
        RECT 0.625 1.720 3.225 1.890 ;
        RECT 3.395 1.820 3.725 2.905 ;
        RECT 0.625 1.630 0.795 1.720 ;
        RECT 0.425 1.300 0.795 1.630 ;
        RECT 0.625 1.020 0.795 1.300 ;
        RECT 0.625 0.850 2.880 1.020 ;
        RECT 0.650 0.085 1.050 0.680 ;
        RECT 2.200 0.430 2.880 0.850 ;
        RECT 3.370 0.085 3.700 1.040 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a32o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a32o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a32o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 2.915 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.015 1.350 2.345 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.445 1.350 1.775 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.350 3.715 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.300 4.215 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.290 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.550600 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.820 0.935 2.150 ;
        RECT 0.725 1.150 0.935 1.820 ;
        RECT 0.615 0.330 0.935 1.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.660 0.445 3.245 ;
        RECT 1.100 2.660 1.510 3.245 ;
        RECT 0.225 2.320 1.275 2.490 ;
        RECT 0.225 1.650 0.395 2.320 ;
        RECT 1.105 2.120 1.275 2.320 ;
        RECT 1.715 2.460 2.045 2.860 ;
        RECT 2.265 2.630 2.645 3.245 ;
        RECT 2.875 2.905 4.205 3.075 ;
        RECT 2.875 2.460 3.205 2.905 ;
        RECT 1.715 2.290 3.205 2.460 ;
        RECT 3.375 2.120 3.705 2.735 ;
        RECT 1.105 1.950 3.705 2.120 ;
        RECT 3.875 1.950 4.205 2.905 ;
        RECT 0.225 1.320 0.555 1.650 ;
        RECT 1.105 1.180 1.275 1.950 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 1.105 1.010 3.105 1.180 ;
        RECT 1.185 0.085 1.515 0.840 ;
        RECT 2.775 0.350 3.105 1.010 ;
        RECT 3.850 0.085 4.180 1.130 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a32o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a32o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.635 1.450 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.180 1.950 6.595 2.120 ;
        RECT 5.180 1.790 5.350 1.950 ;
        RECT 4.440 1.470 5.350 1.790 ;
        RECT 6.425 1.770 6.595 1.950 ;
        RECT 6.425 1.440 6.825 1.770 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 7.065 1.450 8.035 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.450 3.715 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.450 2.835 1.780 ;
        RECT 2.570 0.425 2.740 1.450 ;
        RECT 4.085 0.425 4.415 0.585 ;
        RECT 2.570 0.255 4.415 0.425 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.310 1.380 4.685 1.465 ;
        RECT 3.310 1.320 8.155 1.380 ;
        RECT 0.005 0.245 8.155 1.320 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.780 8.350 3.520 ;
        RECT -0.190 1.660 3.100 1.780 ;
        RECT 4.895 1.660 8.350 1.780 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.097500 ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.020 0.815 2.980 ;
        RECT 1.515 2.020 1.795 3.000 ;
        RECT 0.565 1.850 1.795 2.020 ;
        RECT 0.565 1.650 0.815 1.850 ;
        RECT 0.125 1.480 0.815 1.650 ;
        RECT 0.125 1.180 0.355 1.480 ;
        RECT 0.125 0.930 1.900 1.180 ;
        RECT 0.615 0.410 0.820 0.930 ;
        RECT 1.570 0.430 1.900 0.930 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.015 2.190 1.345 3.245 ;
        RECT 1.965 2.290 2.295 3.245 ;
        RECT 2.525 2.905 4.925 3.075 ;
        RECT 2.525 2.290 2.855 2.905 ;
        RECT 3.025 2.120 3.355 2.735 ;
        RECT 3.525 2.290 3.855 2.905 ;
        RECT 4.025 2.120 4.355 2.735 ;
        RECT 2.015 1.950 4.355 2.120 ;
        RECT 4.595 2.460 4.925 2.905 ;
        RECT 5.210 2.630 5.615 3.245 ;
        RECT 5.785 2.460 6.115 2.900 ;
        RECT 6.285 2.630 6.645 3.245 ;
        RECT 6.815 2.460 7.095 3.000 ;
        RECT 4.595 2.290 7.095 2.460 ;
        RECT 7.265 2.290 7.545 3.245 ;
        RECT 4.595 1.960 4.925 2.290 ;
        RECT 6.765 2.120 7.095 2.290 ;
        RECT 7.715 2.120 8.045 2.980 ;
        RECT 6.765 1.950 8.045 2.120 ;
        RECT 2.015 1.680 2.185 1.950 ;
        RECT 0.985 1.350 2.185 1.680 ;
        RECT 3.885 1.280 4.055 1.950 ;
        RECT 0.115 0.085 0.445 0.760 ;
        RECT 0.990 0.085 1.400 0.760 ;
        RECT 2.070 0.085 2.400 1.180 ;
        RECT 2.910 0.925 3.240 1.210 ;
        RECT 3.420 1.110 6.130 1.280 ;
        RECT 3.420 1.095 3.750 1.110 ;
        RECT 2.910 0.755 4.180 0.925 ;
        RECT 4.350 0.755 4.755 0.940 ;
        RECT 2.910 0.595 3.240 0.755 ;
        RECT 4.585 0.085 4.755 0.755 ;
        RECT 4.940 0.425 5.190 0.940 ;
        RECT 5.370 0.765 5.620 0.940 ;
        RECT 5.800 0.935 6.130 1.110 ;
        RECT 6.310 0.765 6.560 1.270 ;
        RECT 5.370 0.595 6.560 0.765 ;
        RECT 6.740 1.100 8.045 1.270 ;
        RECT 6.740 0.425 6.990 1.100 ;
        RECT 4.940 0.255 6.990 0.425 ;
        RECT 7.190 0.085 7.545 0.920 ;
        RECT 7.715 0.590 8.045 1.100 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__a32o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a32oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a32oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.180 1.855 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.440 2.525 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.765 1.180 3.235 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.180 1.315 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.180 0.445 1.550 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.330 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.998800 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.890 0.945 2.735 ;
        RECT 1.590 1.890 2.275 2.150 ;
        RECT 0.615 1.720 2.275 1.890 ;
        RECT 0.615 1.010 0.785 1.720 ;
        RECT 0.615 0.350 1.830 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.905 1.445 3.075 ;
        RECT 0.115 1.820 0.445 2.905 ;
        RECT 1.115 2.490 1.445 2.905 ;
        RECT 1.675 2.660 2.345 3.245 ;
        RECT 2.515 2.490 2.795 2.980 ;
        RECT 1.115 2.320 2.795 2.490 ;
        RECT 1.115 2.060 1.420 2.320 ;
        RECT 2.465 1.820 2.795 2.320 ;
        RECT 2.995 1.820 3.245 3.245 ;
        RECT 0.115 0.085 0.445 1.010 ;
        RECT 2.890 0.085 3.220 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a32oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a32oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.180 2.775 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.375 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 5.785 1.180 6.115 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.180 2.275 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.630 0.355 1.780 ;
        RECT 0.125 1.300 1.090 1.630 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 6.235 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.192800 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.970 0.945 2.735 ;
        RECT 1.615 1.970 1.945 2.735 ;
        RECT 0.615 1.890 1.945 1.970 ;
        RECT 0.615 1.800 3.235 1.890 ;
        RECT 1.615 1.720 3.235 1.800 ;
        RECT 3.005 1.235 3.235 1.720 ;
        RECT 3.005 1.010 3.205 1.235 ;
        RECT 1.455 0.840 3.205 1.010 ;
        RECT 1.455 0.595 1.785 0.840 ;
        RECT 3.015 0.595 3.205 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.115 2.905 2.400 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 1.115 2.140 1.445 2.905 ;
        RECT 2.115 2.230 2.400 2.905 ;
        RECT 2.570 2.400 3.280 3.245 ;
        RECT 3.450 2.230 3.735 2.980 ;
        RECT 3.905 2.290 4.250 3.245 ;
        RECT 2.115 2.120 3.735 2.230 ;
        RECT 4.420 2.120 4.875 2.980 ;
        RECT 2.115 2.060 4.875 2.120 ;
        RECT 5.045 2.060 5.375 3.245 ;
        RECT 3.405 1.950 4.875 2.060 ;
        RECT 4.545 1.890 4.875 1.950 ;
        RECT 5.545 1.890 5.875 2.980 ;
        RECT 4.545 1.720 5.875 1.890 ;
        RECT 0.115 0.960 1.275 1.130 ;
        RECT 0.115 0.350 0.365 0.960 ;
        RECT 0.545 0.085 0.875 0.790 ;
        RECT 1.105 0.425 1.275 0.960 ;
        RECT 1.955 0.425 2.285 0.670 ;
        RECT 1.105 0.255 2.285 0.425 ;
        RECT 2.515 0.425 2.845 0.670 ;
        RECT 3.375 0.425 3.705 1.130 ;
        RECT 3.875 1.010 5.615 1.180 ;
        RECT 3.875 0.595 4.205 1.010 ;
        RECT 4.375 0.425 4.705 0.840 ;
        RECT 2.515 0.255 4.705 0.425 ;
        RECT 4.935 0.085 5.185 0.840 ;
        RECT 5.365 0.350 5.615 1.010 ;
        RECT 5.795 0.085 6.125 1.010 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__a32oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a32oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a32oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 5.805 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.735 1.350 8.515 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.350 10.435 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 4.195 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.795 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.560 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 10.555 1.240 ;
        RECT 0.000 0.000 10.560 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.750 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.560 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.387000 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 0.945 2.735 ;
        RECT 1.515 2.120 1.845 2.735 ;
        RECT 2.515 2.120 2.845 2.735 ;
        RECT 3.515 2.120 3.845 2.735 ;
        RECT 0.615 1.950 6.350 2.120 ;
        RECT 2.400 1.130 5.150 1.180 ;
        RECT 6.180 1.130 6.350 1.950 ;
        RECT 2.400 1.010 6.350 1.130 ;
        RECT 2.400 0.880 3.660 1.010 ;
        RECT 2.400 0.595 2.730 0.880 ;
        RECT 4.820 0.770 6.350 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.560 3.415 ;
        RECT 0.115 2.905 4.345 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 1.145 2.290 1.315 2.905 ;
        RECT 2.015 2.290 2.345 2.905 ;
        RECT 3.015 2.290 3.345 2.905 ;
        RECT 4.015 2.460 4.345 2.905 ;
        RECT 4.605 2.630 4.935 3.245 ;
        RECT 5.105 2.460 5.435 2.980 ;
        RECT 5.605 2.630 5.935 3.245 ;
        RECT 6.105 2.460 6.435 2.980 ;
        RECT 6.605 2.630 6.935 3.245 ;
        RECT 7.105 2.460 7.435 2.980 ;
        RECT 4.015 2.290 7.435 2.460 ;
        RECT 7.605 2.290 7.935 3.245 ;
        RECT 7.105 2.120 7.435 2.290 ;
        RECT 8.105 2.120 8.435 2.980 ;
        RECT 8.605 2.290 8.935 3.245 ;
        RECT 9.105 2.120 9.435 2.980 ;
        RECT 9.605 2.290 9.935 3.245 ;
        RECT 10.110 2.120 10.440 2.980 ;
        RECT 7.105 1.950 10.440 2.120 ;
        RECT 0.115 1.010 2.220 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.125 0.350 1.295 1.010 ;
        RECT 1.475 0.085 1.805 0.840 ;
        RECT 2.050 0.425 2.220 1.010 ;
        RECT 6.540 1.010 9.935 1.180 ;
        RECT 6.540 0.850 7.735 1.010 ;
        RECT 2.900 0.425 3.230 0.710 ;
        RECT 3.760 0.425 4.090 0.710 ;
        RECT 2.050 0.255 4.090 0.425 ;
        RECT 4.320 0.600 4.650 0.840 ;
        RECT 6.540 0.770 6.870 0.850 ;
        RECT 7.835 0.600 8.165 0.680 ;
        RECT 4.320 0.350 8.165 0.600 ;
        RECT 8.395 0.085 8.725 0.840 ;
        RECT 8.905 0.350 9.075 1.010 ;
        RECT 9.255 0.085 9.585 0.840 ;
        RECT 9.765 0.350 9.935 1.010 ;
        RECT 10.115 0.085 10.445 1.130 ;
        RECT 0.000 -0.085 10.560 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
  END
END sky130_fd_sc_hs__a32oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a41o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a41o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.450 2.355 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.440 2.895 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.135 1.180 3.715 1.550 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.180 4.215 1.550 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.450 1.815 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.270 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.040800 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.820 0.445 2.980 ;
        RECT 0.115 0.940 0.355 1.820 ;
        RECT 0.115 0.290 1.120 0.940 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.645 1.820 0.895 3.245 ;
        RECT 1.145 1.950 1.635 2.980 ;
        RECT 1.805 2.120 2.135 2.980 ;
        RECT 2.305 2.290 2.635 3.245 ;
        RECT 2.835 2.120 3.165 2.980 ;
        RECT 1.805 1.950 3.165 2.120 ;
        RECT 3.335 2.060 3.665 3.245 ;
        RECT 1.145 1.550 1.315 1.950 ;
        RECT 2.835 1.890 3.165 1.950 ;
        RECT 3.855 1.890 4.185 2.980 ;
        RECT 2.835 1.720 4.185 1.890 ;
        RECT 0.575 1.280 1.315 1.550 ;
        RECT 0.575 1.110 2.120 1.280 ;
        RECT 1.290 0.085 1.620 0.940 ;
        RECT 1.790 0.350 2.120 1.110 ;
        RECT 3.830 0.085 4.160 1.010 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a41o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a41o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a41o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.450 2.355 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.440 1.815 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.845 0.440 1.315 1.550 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.455 1.550 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.450 2.925 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.639400 ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.820 4.185 2.980 ;
        RECT 4.015 0.940 4.185 1.820 ;
        RECT 3.385 0.770 4.185 0.940 ;
        RECT 3.385 0.350 3.715 0.770 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 1.890 0.445 2.980 ;
        RECT 0.615 2.060 0.945 3.245 ;
        RECT 1.115 2.120 1.445 2.980 ;
        RECT 1.615 2.290 2.125 3.245 ;
        RECT 2.295 2.120 2.625 2.980 ;
        RECT 1.115 1.950 2.625 2.120 ;
        RECT 2.795 2.120 3.125 2.980 ;
        RECT 3.355 2.270 3.685 3.245 ;
        RECT 2.795 1.950 3.265 2.120 ;
        RECT 1.115 1.890 1.445 1.950 ;
        RECT 0.115 1.720 1.445 1.890 ;
        RECT 3.095 1.550 3.265 1.950 ;
        RECT 4.355 1.820 4.685 3.245 ;
        RECT 3.095 1.280 3.845 1.550 ;
        RECT 2.230 1.110 3.845 1.280 ;
        RECT 0.150 0.085 0.480 1.010 ;
        RECT 2.230 0.350 2.560 1.110 ;
        RECT 2.790 0.085 3.120 0.940 ;
        RECT 3.885 0.085 4.685 0.600 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__a41o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a41o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a41o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.450 4.195 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 4.900 1.450 5.635 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.450 7.075 1.780 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 7.325 1.450 8.035 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.550 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 3.495 1.360 ;
        RECT 0.005 0.245 8.155 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.840 3.305 2.120 ;
        RECT 2.555 1.170 3.305 1.840 ;
        RECT 1.550 1.000 3.305 1.170 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 2.905 1.395 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 0.615 1.950 0.890 2.735 ;
        RECT 0.720 1.670 0.890 1.950 ;
        RECT 1.065 2.460 1.395 2.905 ;
        RECT 1.625 2.630 1.955 3.245 ;
        RECT 2.525 2.630 2.855 3.245 ;
        RECT 3.425 2.650 3.775 3.245 ;
        RECT 4.045 2.460 4.375 2.980 ;
        RECT 1.065 2.290 4.375 2.460 ;
        RECT 4.635 2.290 5.095 3.245 ;
        RECT 1.065 1.940 1.395 2.290 ;
        RECT 4.045 2.120 4.375 2.290 ;
        RECT 5.265 2.120 5.595 2.980 ;
        RECT 5.765 2.290 6.095 3.245 ;
        RECT 6.265 2.120 6.595 2.980 ;
        RECT 6.765 2.290 7.095 3.245 ;
        RECT 7.265 2.120 7.595 2.980 ;
        RECT 4.045 1.950 7.595 2.120 ;
        RECT 7.795 1.950 8.045 3.245 ;
        RECT 0.720 1.340 2.385 1.670 ;
        RECT 0.720 1.250 1.225 1.340 ;
        RECT 0.110 0.085 0.360 1.250 ;
        RECT 0.540 0.830 1.225 1.250 ;
        RECT 0.540 0.660 3.645 0.830 ;
        RECT 3.815 0.770 4.845 1.150 ;
        RECT 5.025 1.110 6.680 1.280 ;
        RECT 5.025 0.770 5.285 1.110 ;
        RECT 3.815 0.700 3.985 0.770 ;
        RECT 0.540 0.470 0.870 0.660 ;
        RECT 1.045 0.085 1.375 0.490 ;
        RECT 2.055 0.085 2.385 0.490 ;
        RECT 3.055 0.085 3.305 0.490 ;
        RECT 3.475 0.425 3.645 0.660 ;
        RECT 4.675 0.600 4.845 0.770 ;
        RECT 5.455 0.600 5.785 0.940 ;
        RECT 4.165 0.425 4.495 0.600 ;
        RECT 3.475 0.255 4.495 0.425 ;
        RECT 4.675 0.330 5.785 0.600 ;
        RECT 6.000 0.425 6.330 0.940 ;
        RECT 6.510 0.595 6.680 1.110 ;
        RECT 6.860 1.110 8.050 1.280 ;
        RECT 6.860 0.425 7.110 1.110 ;
        RECT 6.000 0.255 7.110 0.425 ;
        RECT 7.290 0.085 7.620 0.940 ;
        RECT 7.790 0.350 8.050 1.110 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__a41o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a41oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a41oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.300 3.255 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.195 1.350 2.755 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 1.955 1.780 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.350 1.335 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.330 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.752200 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.115 1.950 0.835 2.120 ;
        RECT 0.605 1.130 0.835 1.950 ;
        RECT 0.115 0.960 3.220 1.130 ;
        RECT 0.115 0.350 0.445 0.960 ;
        RECT 2.890 0.350 3.220 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.615 2.460 0.945 2.980 ;
        RECT 1.115 2.630 1.785 3.245 ;
        RECT 1.445 2.460 1.785 2.630 ;
        RECT 2.405 2.460 2.745 3.245 ;
        RECT 0.615 2.290 1.275 2.460 ;
        RECT 2.915 2.290 3.245 2.980 ;
        RECT 1.105 1.950 3.245 2.290 ;
        RECT 0.615 0.085 1.260 0.680 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a41oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a41oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a41oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.430 1.795 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.630 3.715 1.780 ;
        RECT 2.665 1.300 3.715 1.630 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 4.675 1.780 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.350 5.635 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.085 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 1.055 1.290 ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.810100 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 0.945 2.735 ;
        RECT 0.615 1.950 2.135 2.120 ;
        RECT 1.965 1.650 2.135 1.950 ;
        RECT 1.965 1.260 2.275 1.650 ;
        RECT 1.685 1.180 2.275 1.260 ;
        RECT 0.615 1.090 2.275 1.180 ;
        RECT 0.615 1.010 1.935 1.090 ;
        RECT 0.615 0.400 0.945 1.010 ;
        RECT 1.685 0.595 1.935 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 2.905 1.445 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 1.115 2.460 1.445 2.905 ;
        RECT 1.615 2.650 2.135 3.245 ;
        RECT 2.305 2.460 2.635 2.980 ;
        RECT 1.115 2.290 2.635 2.460 ;
        RECT 2.805 2.290 3.135 3.245 ;
        RECT 2.305 2.120 2.635 2.290 ;
        RECT 3.305 2.120 3.635 2.980 ;
        RECT 3.805 2.290 4.135 3.245 ;
        RECT 4.305 2.120 4.670 3.000 ;
        RECT 4.840 2.290 5.170 3.245 ;
        RECT 5.340 2.120 5.645 3.000 ;
        RECT 2.305 1.950 5.645 2.120 ;
        RECT 2.305 1.820 2.635 1.950 ;
        RECT 0.115 0.085 0.445 1.180 ;
        RECT 4.465 1.130 5.645 1.180 ;
        RECT 2.965 0.920 3.295 1.080 ;
        RECT 1.175 0.425 1.505 0.840 ;
        RECT 2.105 0.750 3.295 0.920 ;
        RECT 3.525 1.010 5.645 1.130 ;
        RECT 3.525 0.850 4.635 1.010 ;
        RECT 2.105 0.425 2.355 0.750 ;
        RECT 3.955 0.580 4.285 0.680 ;
        RECT 1.175 0.255 2.355 0.425 ;
        RECT 2.535 0.330 4.285 0.580 ;
        RECT 4.465 0.350 4.635 0.850 ;
        RECT 4.815 0.085 5.145 0.840 ;
        RECT 5.315 0.350 5.645 1.010 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__a41oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a41oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a41oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.285 1.350 3.295 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.650 4.675 1.780 ;
        RECT 3.965 1.320 5.620 1.650 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.350 8.035 1.780 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.350 9.955 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.430 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 10.075 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.447600 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 0.945 2.735 ;
        RECT 1.645 2.120 1.815 2.735 ;
        RECT 0.615 1.950 3.715 2.120 ;
        RECT 1.645 1.820 2.105 1.950 ;
        RECT 1.815 1.180 2.105 1.820 ;
        RECT 3.465 1.550 3.715 1.950 ;
        RECT 0.545 1.010 2.435 1.180 ;
        RECT 0.545 0.350 0.875 1.010 ;
        RECT 2.105 0.595 2.435 1.010 ;
        RECT 3.465 1.000 3.635 1.550 ;
        RECT 3.305 0.595 3.635 1.000 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.115 2.905 2.345 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 1.115 2.290 1.445 2.905 ;
        RECT 2.015 2.460 2.345 2.905 ;
        RECT 2.515 2.630 2.845 3.245 ;
        RECT 3.015 2.460 3.345 2.980 ;
        RECT 3.545 2.630 3.795 3.245 ;
        RECT 3.970 2.460 4.300 2.980 ;
        RECT 2.015 2.290 4.300 2.460 ;
        RECT 4.500 2.290 4.750 3.245 ;
        RECT 3.970 2.120 4.300 2.290 ;
        RECT 4.930 2.120 5.260 2.980 ;
        RECT 5.460 2.290 5.710 3.245 ;
        RECT 5.880 2.120 6.210 2.980 ;
        RECT 6.410 2.290 6.660 3.245 ;
        RECT 6.830 2.120 7.160 2.980 ;
        RECT 7.360 2.290 7.610 3.245 ;
        RECT 7.780 2.120 8.110 2.980 ;
        RECT 8.280 2.290 8.530 3.245 ;
        RECT 8.730 2.120 9.060 2.980 ;
        RECT 9.260 2.290 9.430 3.245 ;
        RECT 9.630 2.120 9.960 2.980 ;
        RECT 3.970 1.950 9.960 2.120 ;
        RECT 4.930 1.820 5.260 1.950 ;
        RECT 0.115 0.085 0.365 1.130 ;
        RECT 1.045 0.085 1.375 0.840 ;
        RECT 1.605 0.425 1.935 0.840 ;
        RECT 2.605 0.425 3.135 1.130 ;
        RECT 3.805 0.620 4.135 1.130 ;
        RECT 4.305 0.790 7.775 1.130 ;
        RECT 7.445 0.770 7.775 0.790 ;
        RECT 7.955 1.010 9.965 1.180 ;
        RECT 3.805 0.425 5.925 0.620 ;
        RECT 1.605 0.255 5.925 0.425 ;
        RECT 6.155 0.600 6.485 0.620 ;
        RECT 7.955 0.600 8.125 1.010 ;
        RECT 6.155 0.350 8.125 0.600 ;
        RECT 8.305 0.085 8.635 0.840 ;
        RECT 8.815 0.350 8.985 1.010 ;
        RECT 9.165 0.085 9.495 0.840 ;
        RECT 9.715 0.350 9.965 1.010 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__a41oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a211o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a211o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.450 2.755 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.450 1.835 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.570 2.275 0.670 ;
        RECT 2.045 0.255 2.875 0.570 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.385 0.255 3.715 0.670 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.300 1.240 3.630 1.450 ;
        RECT 0.735 0.245 3.630 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.435 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.435 1.075 1.130 ;
        RECT 0.825 0.345 1.075 0.435 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.635 1.820 0.885 3.245 ;
        RECT 1.355 2.120 1.685 2.980 ;
        RECT 1.885 2.290 2.085 3.245 ;
        RECT 2.285 2.120 2.615 2.980 ;
        RECT 1.355 1.950 2.615 2.120 ;
        RECT 0.425 1.400 1.415 1.650 ;
        RECT 1.245 1.280 1.415 1.400 ;
        RECT 3.125 1.280 3.540 2.980 ;
        RECT 1.245 1.110 3.540 1.280 ;
        RECT 2.280 1.080 3.540 1.110 ;
        RECT 1.255 0.085 1.705 0.940 ;
        RECT 2.280 0.840 2.610 1.080 ;
        RECT 2.780 0.740 3.215 0.910 ;
        RECT 3.045 0.085 3.215 0.740 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a211o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a211o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a211o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.260 2.535 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.260 1.875 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.745 1.260 3.235 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.450 3.735 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 0.245 3.830 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.180 0.835 2.980 ;
        RECT 0.575 1.010 0.980 1.180 ;
        RECT 0.810 0.350 0.980 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.125 1.820 0.375 3.245 ;
        RECT 1.025 2.290 1.355 3.245 ;
        RECT 1.545 2.460 1.875 2.980 ;
        RECT 2.075 2.630 2.365 3.245 ;
        RECT 2.535 2.460 2.865 2.980 ;
        RECT 1.545 2.290 2.865 2.460 ;
        RECT 3.405 2.120 3.735 2.980 ;
        RECT 1.165 1.950 3.735 2.120 ;
        RECT 1.165 1.680 1.335 1.950 ;
        RECT 1.005 1.350 1.335 1.680 ;
        RECT 1.165 1.090 1.335 1.350 ;
        RECT 3.490 1.090 3.740 1.130 ;
        RECT 1.165 0.920 3.740 1.090 ;
        RECT 0.300 0.085 0.630 0.840 ;
        RECT 1.160 0.350 1.870 0.750 ;
        RECT 2.330 0.350 2.700 0.920 ;
        RECT 2.870 0.350 3.310 0.750 ;
        RECT 3.490 0.350 3.740 0.920 ;
        RECT 1.160 0.085 1.330 0.350 ;
        RECT 2.870 0.085 3.040 0.350 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a211o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a211o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.450 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 0.505 5.125 0.670 ;
        RECT 4.925 0.255 5.320 0.505 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.995 1.890 4.195 2.150 ;
        RECT 2.785 1.720 4.515 1.890 ;
        RECT 2.785 1.470 3.105 1.720 ;
        RECT 3.965 1.470 4.515 1.720 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.450 1.210 3.780 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.920 1.310 7.005 1.385 ;
        RECT 3.445 1.240 7.005 1.310 ;
        RECT 0.730 0.245 7.005 1.240 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.675 1.890 0.925 2.980 ;
        RECT 1.575 1.890 1.905 2.980 ;
        RECT 0.675 1.720 1.905 1.890 ;
        RECT 0.675 1.410 0.925 1.720 ;
        RECT 0.675 1.240 1.795 1.410 ;
        RECT 1.330 0.960 1.795 1.240 ;
        RECT 1.330 0.790 2.370 0.960 ;
        RECT 1.330 0.350 1.500 0.790 ;
        RECT 2.180 0.545 2.370 0.790 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.225 1.820 0.475 3.245 ;
        RECT 1.125 2.060 1.375 3.245 ;
        RECT 2.105 1.820 2.275 3.245 ;
        RECT 2.545 2.570 2.875 2.780 ;
        RECT 3.045 2.740 4.300 2.990 ;
        RECT 4.500 2.570 4.710 2.990 ;
        RECT 2.545 2.400 4.710 2.570 ;
        RECT 4.880 2.400 5.555 3.245 ;
        RECT 4.420 2.230 4.710 2.400 ;
        RECT 5.725 2.230 5.960 2.980 ;
        RECT 6.130 2.290 6.460 3.245 ;
        RECT 2.445 2.060 3.825 2.230 ;
        RECT 4.420 2.120 5.960 2.230 ;
        RECT 6.630 2.120 6.910 2.980 ;
        RECT 4.420 2.060 6.910 2.120 ;
        RECT 2.445 1.550 2.615 2.060 ;
        RECT 5.680 1.950 6.910 2.060 ;
        RECT 6.580 1.940 6.910 1.950 ;
        RECT 1.965 1.300 2.615 1.550 ;
        RECT 1.965 1.130 3.280 1.300 ;
        RECT 0.820 0.085 1.150 1.050 ;
        RECT 3.040 1.040 3.280 1.130 ;
        RECT 3.960 1.110 6.055 1.280 ;
        RECT 3.960 1.040 4.245 1.110 ;
        RECT 1.680 0.085 2.010 0.620 ;
        RECT 2.540 0.085 2.870 0.960 ;
        RECT 3.040 0.870 4.245 1.040 ;
        RECT 5.725 1.015 6.055 1.110 ;
        RECT 3.040 0.450 3.280 0.870 ;
        RECT 3.460 0.085 3.790 0.700 ;
        RECT 3.960 0.595 4.245 0.870 ;
        RECT 4.425 0.085 4.755 0.940 ;
        RECT 6.235 0.845 6.405 1.275 ;
        RECT 5.295 0.675 6.405 0.845 ;
        RECT 6.235 0.595 6.405 0.675 ;
        RECT 6.585 0.085 6.915 1.275 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__a211o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a211oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a211oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.350 1.335 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.465 1.350 0.835 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.180 2.775 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.250 0.245 2.630 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.792700 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.820 2.565 2.980 ;
        RECT 2.045 1.180 2.215 1.820 ;
        RECT 1.085 1.025 2.215 1.180 ;
        RECT 1.085 1.010 2.275 1.025 ;
        RECT 1.085 0.810 2.540 1.010 ;
        RECT 1.085 0.350 1.500 0.810 ;
        RECT 2.210 0.350 2.540 0.810 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.315 2.120 0.645 2.980 ;
        RECT 0.815 2.290 1.135 3.245 ;
        RECT 1.305 2.120 1.635 2.980 ;
        RECT 0.315 1.950 1.635 2.120 ;
        RECT 0.340 0.085 0.670 1.130 ;
        RECT 1.670 0.085 2.040 0.640 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__a211oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a211oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a211oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.480 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.430 2.275 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.180 3.715 1.550 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.180 4.675 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.245 4.200 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.076000 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.890 4.145 2.735 ;
        RECT 2.525 1.720 4.145 1.890 ;
        RECT 2.525 1.260 2.755 1.720 ;
        RECT 0.650 1.090 2.755 1.260 ;
        RECT 0.650 0.635 0.830 1.090 ;
        RECT 2.585 1.010 2.755 1.090 ;
        RECT 2.585 0.840 3.590 1.010 ;
        RECT 2.960 0.330 3.590 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.105 1.820 0.355 3.245 ;
        RECT 0.555 2.120 0.805 2.980 ;
        RECT 1.005 2.290 1.335 3.245 ;
        RECT 1.535 2.230 1.705 2.980 ;
        RECT 1.905 2.400 2.235 3.245 ;
        RECT 2.465 2.905 4.595 3.075 ;
        RECT 2.465 2.400 2.795 2.905 ;
        RECT 2.965 2.230 3.245 2.735 ;
        RECT 1.535 2.120 3.245 2.230 ;
        RECT 0.555 2.060 3.245 2.120 ;
        RECT 3.445 2.060 3.615 2.905 ;
        RECT 0.555 1.950 2.355 2.060 ;
        RECT 0.555 1.820 0.805 1.950 ;
        RECT 4.345 1.820 4.595 2.905 ;
        RECT 0.150 0.425 0.480 1.010 ;
        RECT 1.010 0.750 2.240 0.920 ;
        RECT 1.010 0.425 1.260 0.750 ;
        RECT 0.150 0.255 1.260 0.425 ;
        RECT 1.440 0.330 1.810 0.580 ;
        RECT 1.990 0.330 2.240 0.750 ;
        RECT 1.440 0.085 1.610 0.330 ;
        RECT 2.460 0.085 2.790 0.670 ;
        RECT 3.760 0.085 4.090 1.010 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__a211oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a211oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.350 3.855 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 2.275 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.300 6.115 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.350 7.555 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.330 0.245 4.300 1.240 ;
        RECT 5.290 0.245 7.520 1.240 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.685800 ;
    PORT
      LAYER li1 ;
        RECT 6.795 2.120 6.965 2.735 ;
        RECT 7.695 2.120 7.895 2.735 ;
        RECT 6.795 1.950 7.895 2.120 ;
        RECT 7.725 1.180 8.515 1.950 ;
        RECT 6.320 1.130 8.515 1.180 ;
        RECT 2.570 1.010 8.515 1.130 ;
        RECT 2.570 0.960 6.490 1.010 ;
        RECT 2.570 0.785 3.760 0.960 ;
        RECT 5.380 0.350 5.630 0.960 ;
        RECT 6.320 0.350 6.490 0.960 ;
        RECT 7.180 0.350 8.515 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.345 2.120 0.675 2.980 ;
        RECT 0.875 2.290 1.045 3.245 ;
        RECT 1.245 2.120 1.495 2.980 ;
        RECT 1.695 2.290 2.025 3.245 ;
        RECT 2.225 2.120 2.395 2.980 ;
        RECT 2.595 2.290 2.925 3.245 ;
        RECT 3.125 2.120 3.295 2.980 ;
        RECT 3.495 2.290 3.825 3.245 ;
        RECT 4.025 2.120 4.275 2.980 ;
        RECT 4.465 2.905 8.395 3.075 ;
        RECT 4.465 2.290 4.795 2.905 ;
        RECT 4.995 2.120 5.165 2.735 ;
        RECT 5.365 2.290 5.695 2.905 ;
        RECT 5.895 2.120 6.145 2.735 ;
        RECT 0.345 1.950 6.145 2.120 ;
        RECT 6.315 1.950 6.595 2.905 ;
        RECT 7.165 2.290 7.495 2.905 ;
        RECT 8.065 2.120 8.395 2.905 ;
        RECT 4.025 1.820 4.275 1.950 ;
        RECT 0.420 1.010 2.390 1.180 ;
        RECT 0.420 0.350 0.670 1.010 ;
        RECT 0.850 0.085 1.180 0.840 ;
        RECT 1.360 0.350 1.530 1.010 ;
        RECT 1.710 0.085 2.040 0.840 ;
        RECT 2.220 0.615 2.390 1.010 ;
        RECT 2.220 0.350 4.190 0.615 ;
        RECT 5.810 0.085 6.140 0.790 ;
        RECT 6.670 0.085 7.000 0.840 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__a211oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a221o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a221o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.470 2.295 1.800 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.375 1.350 1.795 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.455 2.985 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.195 1.455 3.715 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.865 0.255 4.195 0.670 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.525 1.165 1.450 1.240 ;
        RECT 3.355 1.165 4.280 1.385 ;
        RECT 0.525 0.245 4.280 1.165 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.820 0.900 2.980 ;
        RECT 0.125 1.130 0.500 1.820 ;
        RECT 0.125 0.350 0.865 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 1.100 1.950 1.350 3.245 ;
        RECT 1.535 2.140 1.785 2.980 ;
        RECT 1.985 2.310 2.315 3.245 ;
        RECT 2.505 2.905 3.685 3.075 ;
        RECT 2.505 2.310 2.785 2.905 ;
        RECT 2.955 2.140 3.285 2.735 ;
        RECT 1.535 1.970 3.285 2.140 ;
        RECT 1.535 1.950 1.785 1.970 ;
        RECT 2.955 1.950 3.285 1.970 ;
        RECT 3.485 1.950 3.685 2.905 ;
        RECT 0.740 1.300 1.205 1.630 ;
        RECT 1.035 1.180 1.205 1.300 ;
        RECT 3.885 1.285 4.215 2.980 ;
        RECT 2.465 1.180 4.215 1.285 ;
        RECT 1.035 1.115 4.215 1.180 ;
        RECT 1.035 1.010 2.860 1.115 ;
        RECT 1.045 0.085 1.965 0.840 ;
        RECT 2.420 0.375 2.860 1.010 ;
        RECT 3.320 0.085 3.690 0.945 ;
        RECT 3.860 0.840 4.215 1.115 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a221o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a221o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a221o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.450 2.275 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.365 1.260 1.765 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.455 1.450 2.760 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.270 1.180 3.695 1.550 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.865 1.180 4.195 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.085 0.245 4.310 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.600 1.970 0.930 2.980 ;
        RECT 0.100 1.800 0.930 1.970 ;
        RECT 0.100 1.130 0.335 1.800 ;
        RECT 0.100 0.960 0.855 1.130 ;
        RECT 0.605 0.350 0.855 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.150 2.140 0.400 3.245 ;
        RECT 1.130 1.950 1.380 3.245 ;
        RECT 1.565 2.120 1.815 2.980 ;
        RECT 2.015 2.290 2.345 3.245 ;
        RECT 2.535 2.905 3.685 3.075 ;
        RECT 2.535 2.400 2.785 2.905 ;
        RECT 2.985 2.230 3.315 2.735 ;
        RECT 2.540 2.120 3.315 2.230 ;
        RECT 1.565 2.060 3.315 2.120 ;
        RECT 3.515 2.060 3.685 2.905 ;
        RECT 1.565 1.950 2.730 2.060 ;
        RECT 3.885 1.890 4.215 2.980 ;
        RECT 2.930 1.720 4.215 1.890 ;
        RECT 0.525 1.300 1.195 1.630 ;
        RECT 1.025 1.090 1.195 1.300 ;
        RECT 2.930 1.130 3.100 1.720 ;
        RECT 2.020 1.090 3.100 1.130 ;
        RECT 1.025 1.010 3.100 1.090 ;
        RECT 1.025 0.920 4.220 1.010 ;
        RECT 2.020 0.840 4.220 0.920 ;
        RECT 0.175 0.085 0.425 0.790 ;
        RECT 1.035 0.085 1.560 0.750 ;
        RECT 2.020 0.350 2.890 0.840 ;
        RECT 3.350 0.085 3.720 0.670 ;
        RECT 3.890 0.350 4.220 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a221o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a221o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a221o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.595 0.565 1.765 1.040 ;
        RECT 1.435 0.255 1.765 0.565 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.505 2.755 0.670 ;
        RECT 2.275 0.255 2.755 0.505 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 8.615 1.300 9.495 1.750 ;
        RECT 9.095 1.210 9.495 1.300 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 0.505 7.045 0.670 ;
        RECT 6.470 0.255 7.045 0.505 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.470 5.735 2.150 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.225 1.385 1.595 1.445 ;
        RECT 0.225 1.370 3.345 1.385 ;
        RECT 6.185 1.370 7.555 1.385 ;
        RECT 0.225 1.150 7.555 1.370 ;
        RECT 0.225 0.245 9.035 1.150 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER met1 ;
        RECT 0.095 1.365 0.385 1.410 ;
        RECT 2.975 1.365 3.265 1.410 ;
        RECT 0.095 1.225 3.265 1.365 ;
        RECT 0.095 1.180 0.385 1.225 ;
        RECT 2.975 1.180 3.265 1.225 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.320 2.260 0.650 3.245 ;
        RECT 0.890 2.430 1.220 2.900 ;
        RECT 1.395 2.600 2.065 3.245 ;
        RECT 2.235 2.530 2.565 2.900 ;
        RECT 2.845 2.700 3.175 3.245 ;
        RECT 3.745 2.700 4.075 3.245 ;
        RECT 4.645 2.700 4.975 3.245 ;
        RECT 5.470 2.905 8.830 3.075 ;
        RECT 5.470 2.700 6.700 2.905 ;
        RECT 6.870 2.530 7.150 2.735 ;
        RECT 2.235 2.430 7.150 2.530 ;
        RECT 0.890 2.360 7.150 2.430 ;
        RECT 0.890 2.260 2.565 2.360 ;
        RECT 2.850 2.090 4.525 2.190 ;
        RECT 0.125 1.920 4.525 2.090 ;
        RECT 0.125 1.180 0.355 1.920 ;
        RECT 5.920 1.770 6.250 2.190 ;
        RECT 6.820 2.110 7.150 2.360 ;
        RECT 7.425 2.280 7.755 2.905 ;
        RECT 8.010 2.110 8.380 2.735 ;
        RECT 6.820 1.940 8.380 2.110 ;
        RECT 8.580 1.940 8.830 2.905 ;
        RECT 0.745 1.580 4.880 1.750 ;
        RECT 0.745 1.075 1.075 1.580 ;
        RECT 1.255 1.240 2.760 1.410 ;
        RECT 0.315 0.905 0.565 1.010 ;
        RECT 1.255 0.905 1.425 1.240 ;
        RECT 0.315 0.735 1.425 0.905 ;
        RECT 0.315 0.655 0.565 0.735 ;
        RECT 1.935 0.675 2.330 1.070 ;
        RECT 2.510 0.840 2.760 1.240 ;
        RECT 3.005 1.180 3.235 1.410 ;
        RECT 3.595 1.350 4.880 1.580 ;
        RECT 4.710 1.300 4.880 1.350 ;
        RECT 5.920 1.600 8.445 1.770 ;
        RECT 5.920 1.300 6.090 1.600 ;
        RECT 3.005 1.010 4.540 1.180 ;
        RECT 4.710 1.130 6.090 1.300 ;
        RECT 1.935 0.085 2.105 0.675 ;
        RECT 3.000 0.085 3.250 0.840 ;
        RECT 3.430 0.440 3.760 1.010 ;
        RECT 3.940 0.085 4.110 0.840 ;
        RECT 4.290 0.480 4.540 1.010 ;
        RECT 4.720 0.085 5.440 0.960 ;
        RECT 5.610 0.580 5.940 1.130 ;
        RECT 6.275 0.960 6.525 1.280 ;
        RECT 6.130 0.675 6.525 0.960 ;
        RECT 6.705 1.260 7.935 1.430 ;
        RECT 6.705 0.840 7.035 1.260 ;
        RECT 6.130 0.085 6.300 0.675 ;
        RECT 7.215 0.085 7.465 1.090 ;
        RECT 7.685 0.425 7.935 1.260 ;
        RECT 8.115 0.595 8.445 1.600 ;
        RECT 8.625 0.425 8.925 1.040 ;
        RECT 7.685 0.255 8.925 0.425 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 0.155 1.210 0.325 1.380 ;
        RECT 3.035 1.210 3.205 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
  END
END sky130_fd_sc_hs__a221o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a221oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.350 2.835 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.180 3.715 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.350 2.295 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.350 1.795 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.350 0.875 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.330 0.245 3.590 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.177500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.375 2.980 ;
        RECT 0.125 1.010 2.575 1.180 ;
        RECT 0.125 0.350 1.090 1.010 ;
        RECT 2.160 0.350 2.575 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.575 2.905 2.055 3.075 ;
        RECT 0.575 1.950 0.905 2.905 ;
        RECT 1.275 2.120 1.545 2.735 ;
        RECT 1.725 2.290 2.055 2.905 ;
        RECT 2.255 2.120 2.505 2.980 ;
        RECT 2.675 2.290 3.025 3.245 ;
        RECT 3.195 2.120 3.525 2.980 ;
        RECT 1.275 1.950 3.525 2.120 ;
        RECT 3.195 1.820 3.525 1.950 ;
        RECT 1.260 0.085 1.630 0.825 ;
        RECT 3.170 0.085 3.500 1.010 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a221oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a221oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a221oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.950 5.065 2.120 ;
        RECT 3.405 1.430 3.735 1.950 ;
        RECT 4.895 1.780 5.065 1.950 ;
        RECT 4.895 1.430 5.635 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.430 4.675 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.425 1.950 3.235 2.120 ;
        RECT 1.425 1.680 1.595 1.950 ;
        RECT 1.245 1.430 1.595 1.680 ;
        RECT 2.525 1.550 3.235 1.950 ;
        RECT 2.685 1.430 3.015 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.430 2.275 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.585 1.350 0.915 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.245 5.520 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.172200 ;
    PORT
      LAYER li1 ;
        RECT 0.555 2.120 0.885 2.735 ;
        RECT 0.125 1.950 0.885 2.120 ;
        RECT 0.125 1.180 0.380 1.950 ;
        RECT 1.090 1.180 5.430 1.260 ;
        RECT 0.125 1.090 5.430 1.180 ;
        RECT 0.125 1.010 1.260 1.090 ;
        RECT 0.125 0.350 0.380 1.010 ;
        RECT 1.090 0.350 1.260 1.010 ;
        RECT 2.950 0.350 3.180 1.090 ;
        RECT 5.180 0.350 5.430 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.105 2.980 2.265 3.075 ;
        RECT 0.105 2.905 3.165 2.980 ;
        RECT 0.105 2.290 0.355 2.905 ;
        RECT 1.085 1.850 1.255 2.905 ;
        RECT 1.455 2.460 1.815 2.735 ;
        RECT 2.015 2.630 3.165 2.905 ;
        RECT 3.355 2.630 3.605 3.245 ;
        RECT 3.805 2.460 4.135 2.980 ;
        RECT 4.335 2.630 4.505 3.245 ;
        RECT 4.705 2.460 5.035 2.980 ;
        RECT 1.455 2.290 5.035 2.460 ;
        RECT 5.235 1.950 5.485 3.245 ;
        RECT 0.560 0.085 0.910 0.840 ;
        RECT 1.440 0.750 2.780 0.920 ;
        RECT 1.440 0.350 1.770 0.750 ;
        RECT 1.940 0.085 2.280 0.580 ;
        RECT 2.450 0.330 2.780 0.750 ;
        RECT 3.350 0.750 5.000 0.920 ;
        RECT 3.350 0.330 4.030 0.750 ;
        RECT 4.200 0.085 4.530 0.580 ;
        RECT 4.700 0.330 5.000 0.750 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__a221oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a221oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.430 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.430 4.265 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.430 8.095 1.780 ;
        RECT 6.730 1.350 8.095 1.430 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.350 9.955 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.350 1.875 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.560 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 0.245 10.450 1.240 ;
        RECT 0.000 0.000 10.560 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.750 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.560 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.380200 ;
    PORT
      LAYER li1 ;
        RECT 0.105 2.905 2.235 3.075 ;
        RECT 0.105 1.180 0.355 2.905 ;
        RECT 1.005 2.290 1.335 2.905 ;
        RECT 1.905 2.290 2.235 2.905 ;
        RECT 2.045 1.180 6.530 1.260 ;
        RECT 0.105 1.090 8.210 1.180 ;
        RECT 0.105 1.010 2.295 1.090 ;
        RECT 0.105 0.350 0.495 1.010 ;
        RECT 1.185 0.350 1.355 1.010 ;
        RECT 2.045 0.350 2.295 1.010 ;
        RECT 4.850 0.640 5.040 1.090 ;
        RECT 5.710 0.640 5.900 1.090 ;
        RECT 6.360 0.850 8.210 1.090 ;
        RECT 7.915 0.770 8.210 0.850 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.560 3.415 ;
        RECT 0.555 2.120 0.835 2.735 ;
        RECT 1.505 2.120 1.735 2.735 ;
        RECT 2.615 2.460 2.945 2.980 ;
        RECT 3.145 2.630 3.315 3.245 ;
        RECT 3.515 2.460 3.845 2.980 ;
        RECT 4.045 2.630 4.215 3.245 ;
        RECT 4.415 2.460 4.745 2.980 ;
        RECT 4.945 2.630 5.115 3.245 ;
        RECT 5.315 2.460 5.645 2.980 ;
        RECT 5.815 2.630 6.275 3.245 ;
        RECT 6.445 2.905 10.375 3.075 ;
        RECT 6.445 2.460 6.725 2.905 ;
        RECT 2.615 2.290 6.725 2.460 ;
        RECT 6.895 2.120 7.225 2.735 ;
        RECT 7.395 2.290 7.625 2.905 ;
        RECT 7.795 2.120 8.125 2.735 ;
        RECT 8.295 2.290 8.525 2.905 ;
        RECT 8.695 2.120 9.025 2.735 ;
        RECT 9.195 2.290 9.425 2.905 ;
        RECT 9.595 2.120 9.925 2.735 ;
        RECT 0.555 1.950 9.925 2.120 ;
        RECT 10.125 1.820 10.375 2.905 ;
        RECT 8.390 1.010 10.360 1.180 ;
        RECT 0.675 0.085 1.005 0.840 ;
        RECT 1.535 0.085 1.865 0.840 ;
        RECT 2.630 0.750 4.680 0.920 ;
        RECT 2.630 0.350 2.880 0.750 ;
        RECT 3.060 0.085 3.390 0.580 ;
        RECT 3.570 0.350 3.740 0.750 ;
        RECT 3.920 0.085 4.250 0.580 ;
        RECT 4.430 0.470 4.680 0.750 ;
        RECT 5.210 0.470 5.540 0.920 ;
        RECT 6.070 0.470 6.400 0.680 ;
        RECT 4.430 0.300 6.400 0.470 ;
        RECT 6.590 0.600 6.920 0.680 ;
        RECT 7.450 0.600 7.745 0.680 ;
        RECT 8.390 0.600 8.560 1.010 ;
        RECT 6.590 0.350 8.560 0.600 ;
        RECT 8.740 0.085 9.070 0.840 ;
        RECT 9.250 0.350 9.420 1.010 ;
        RECT 9.600 0.085 9.930 0.840 ;
        RECT 10.110 0.350 10.360 1.010 ;
        RECT 0.000 -0.085 10.560 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
  END
END sky130_fd_sc_hs__a221oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a222o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a222o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.120 3.255 1.520 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.120 3.825 1.545 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.220 1.120 2.755 1.790 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.180 1.930 1.760 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.120 0.550 1.790 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.120 1.390 1.760 ;
    END
  END C2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.850 1.140 4.795 1.240 ;
        RECT 0.030 0.245 4.795 1.140 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 4.355 1.820 4.710 2.980 ;
        RECT 4.540 1.130 4.710 1.820 ;
        RECT 4.355 0.350 4.710 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 2.905 2.590 3.075 ;
        RECT 0.115 1.960 0.445 2.905 ;
        RECT 0.720 1.930 1.050 2.735 ;
        RECT 1.220 1.930 1.550 2.905 ;
        RECT 1.720 2.130 2.050 2.735 ;
        RECT 2.260 2.300 2.590 2.905 ;
        RECT 2.820 2.300 3.150 3.245 ;
        RECT 3.320 2.130 3.650 2.935 ;
        RECT 1.720 1.960 3.650 2.130 ;
        RECT 1.720 1.930 2.050 1.960 ;
        RECT 0.720 0.950 0.890 1.930 ;
        RECT 3.320 1.895 3.650 1.960 ;
        RECT 3.855 1.895 4.185 3.245 ;
        RECT 4.015 1.300 4.370 1.630 ;
        RECT 4.015 0.950 4.185 1.300 ;
        RECT 0.140 0.780 4.185 0.950 ;
        RECT 0.140 0.350 0.470 0.780 ;
        RECT 0.960 0.085 1.805 0.600 ;
        RECT 2.295 0.330 3.130 0.780 ;
        RECT 3.620 0.085 4.185 0.610 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__a222o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a222o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a222o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.350 3.255 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 4.685 1.350 5.155 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.465 1.350 3.795 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 4.445 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.260 1.140 1.780 ;
    END
  END C2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.190 1.180 2.530 1.280 ;
        RECT 0.005 1.140 2.530 1.180 ;
        RECT 0.005 0.245 5.250 1.140 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.695 1.820 2.440 2.200 ;
        RECT 1.695 0.920 2.025 1.820 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.115 2.200 0.365 2.980 ;
        RECT 0.565 2.540 0.895 2.980 ;
        RECT 1.575 2.710 1.905 3.245 ;
        RECT 2.645 2.710 2.975 3.245 ;
        RECT 3.265 2.905 4.665 3.075 ;
        RECT 3.265 2.710 3.630 2.905 ;
        RECT 3.835 2.540 4.165 2.735 ;
        RECT 0.565 2.370 4.165 2.540 ;
        RECT 0.115 1.950 1.525 2.200 ;
        RECT 3.835 1.950 4.165 2.370 ;
        RECT 4.335 1.950 4.665 2.905 ;
        RECT 4.835 1.950 5.165 3.245 ;
        RECT 1.355 1.090 1.525 1.950 ;
        RECT 0.115 0.920 1.525 1.090 ;
        RECT 0.115 0.390 0.365 0.920 ;
        RECT 1.355 0.750 1.525 0.920 ;
        RECT 2.230 1.180 2.560 1.590 ;
        RECT 2.230 1.010 3.750 1.180 ;
        RECT 2.230 0.750 2.400 1.010 ;
        RECT 0.935 0.085 1.185 0.750 ;
        RECT 1.355 0.580 2.400 0.750 ;
        RECT 2.765 0.520 3.095 0.840 ;
        RECT 3.265 0.700 3.750 1.010 ;
        RECT 3.920 1.010 5.140 1.180 ;
        RECT 3.920 0.520 4.090 1.010 ;
        RECT 2.205 0.085 2.535 0.410 ;
        RECT 2.765 0.350 4.090 0.520 ;
        RECT 4.260 0.085 4.590 0.840 ;
        RECT 4.810 0.350 5.140 1.010 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__a222o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a222oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a222oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.120 3.715 1.790 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.180 4.215 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.120 2.875 1.790 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.120 2.305 1.790 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.120 0.595 1.790 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.120 1.315 1.790 ;
    END
  END C2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.245 4.290 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.232000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.130 0.445 2.980 ;
        RECT 1.115 2.130 1.655 2.735 ;
        RECT 0.115 1.960 1.655 2.130 ;
        RECT 1.485 1.780 1.655 1.960 ;
        RECT 1.485 0.950 1.795 1.780 ;
        RECT 0.140 0.780 3.360 0.950 ;
        RECT 0.140 0.350 0.470 0.780 ;
        RECT 2.525 0.330 3.360 0.780 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.615 2.905 2.655 3.075 ;
        RECT 0.615 2.300 0.945 2.905 ;
        RECT 1.825 2.130 2.155 2.735 ;
        RECT 2.325 2.300 2.655 2.905 ;
        RECT 2.825 2.130 3.155 2.980 ;
        RECT 3.325 2.300 3.655 3.245 ;
        RECT 3.875 2.130 4.205 2.980 ;
        RECT 1.825 1.960 4.205 2.130 ;
        RECT 0.960 0.085 2.180 0.600 ;
        RECT 3.850 0.085 4.180 0.950 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a222oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a222oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a222oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.945 1.950 6.055 2.120 ;
        RECT 4.945 1.780 5.115 1.950 ;
        RECT 4.685 1.450 5.115 1.780 ;
        RECT 5.885 1.780 6.055 1.950 ;
        RECT 5.885 1.450 6.455 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.305 1.450 5.635 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.065 1.950 4.275 2.120 ;
        RECT 3.065 1.800 3.235 1.950 ;
        RECT 2.675 1.470 3.235 1.800 ;
        RECT 4.105 1.780 4.275 1.950 ;
        RECT 4.105 1.450 4.475 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.260 3.735 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.165 1.335 1.495 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.665 2.125 1.835 ;
        RECT 0.605 1.495 0.835 1.665 ;
        RECT 0.425 1.165 0.835 1.495 ;
        RECT 1.795 1.130 2.125 1.665 ;
    END
  END C2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 6.690 1.140 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.693200 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.175 0.365 2.980 ;
        RECT 1.065 2.175 1.325 2.735 ;
        RECT 1.995 2.175 2.465 2.735 ;
        RECT 0.085 2.005 2.465 2.175 ;
        RECT 0.085 1.920 0.365 2.005 ;
        RECT 0.085 0.995 0.255 1.920 ;
        RECT 2.295 1.300 2.465 2.005 ;
        RECT 2.295 1.130 2.840 1.300 ;
        RECT 2.510 1.090 2.840 1.130 ;
        RECT 4.450 1.110 6.580 1.280 ;
        RECT 4.450 1.090 4.715 1.110 ;
        RECT 0.085 0.825 1.420 0.995 ;
        RECT 1.090 0.780 1.420 0.825 ;
        RECT 2.510 0.920 4.715 1.090 ;
        RECT 2.510 0.350 2.840 0.920 ;
        RECT 4.450 0.350 4.715 0.920 ;
        RECT 6.320 0.350 6.580 1.110 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.565 2.980 3.335 3.075 ;
        RECT 0.565 2.905 4.325 2.980 ;
        RECT 0.565 2.345 0.895 2.905 ;
        RECT 1.495 2.345 1.825 2.905 ;
        RECT 2.635 2.460 2.805 2.735 ;
        RECT 3.005 2.650 4.325 2.905 ;
        RECT 3.005 2.630 3.335 2.650 ;
        RECT 4.500 2.480 4.715 2.980 ;
        RECT 4.895 2.650 5.255 3.245 ;
        RECT 5.425 2.480 5.655 2.980 ;
        RECT 5.825 2.650 6.155 3.245 ;
        RECT 6.335 2.480 6.605 3.000 ;
        RECT 4.500 2.460 6.605 2.480 ;
        RECT 2.635 2.290 6.605 2.460 ;
        RECT 2.635 1.970 2.805 2.290 ;
        RECT 4.445 1.950 4.775 2.290 ;
        RECT 6.275 1.950 6.605 2.290 ;
        RECT 0.115 0.085 0.480 0.655 ;
        RECT 1.590 0.610 1.780 0.885 ;
        RECT 0.660 0.350 1.780 0.610 ;
        RECT 1.950 0.085 2.280 0.940 ;
        RECT 4.885 0.770 6.150 0.940 ;
        RECT 3.020 0.580 4.270 0.750 ;
        RECT 3.020 0.350 3.270 0.580 ;
        RECT 3.450 0.085 3.840 0.410 ;
        RECT 4.020 0.350 4.270 0.580 ;
        RECT 4.885 0.350 5.215 0.770 ;
        RECT 5.385 0.085 5.715 0.600 ;
        RECT 5.900 0.330 6.150 0.770 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__a222oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a311o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a311o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.440 2.335 0.670 ;
        RECT 2.005 0.255 2.335 0.440 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.450 1.905 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.115 1.450 1.365 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.505 2.725 0.670 ;
        RECT 2.525 0.255 2.875 0.505 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.385 0.255 3.715 0.670 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.265 1.370 3.665 1.385 ;
        RECT 0.265 0.245 3.665 1.370 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.850 0.475 2.980 ;
        RECT 0.125 1.180 0.295 1.850 ;
        RECT 0.125 1.010 0.605 1.180 ;
        RECT 0.355 0.480 0.605 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.645 1.950 1.105 3.245 ;
        RECT 1.275 2.120 1.605 2.980 ;
        RECT 1.805 2.290 2.095 3.245 ;
        RECT 2.265 2.120 2.595 2.980 ;
        RECT 1.275 1.950 2.595 2.120 ;
        RECT 2.265 1.940 2.595 1.950 ;
        RECT 3.105 1.940 3.575 2.980 ;
        RECT 0.480 1.350 0.945 1.680 ;
        RECT 3.245 1.615 3.575 1.940 ;
        RECT 0.775 1.280 0.945 1.350 ;
        RECT 2.240 1.445 3.575 1.615 ;
        RECT 2.240 1.280 2.570 1.445 ;
        RECT 0.775 1.110 2.570 1.280 ;
        RECT 0.785 0.085 1.115 0.940 ;
        RECT 2.240 0.840 2.570 1.110 ;
        RECT 2.750 0.855 3.075 1.185 ;
        RECT 3.245 1.015 3.575 1.445 ;
        RECT 2.895 0.845 3.075 0.855 ;
        RECT 2.895 0.675 3.215 0.845 ;
        RECT 3.045 0.085 3.215 0.675 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__a311o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a311o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a311o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.450 2.835 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.450 2.295 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.260 1.795 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.260 3.715 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.440 4.215 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 0.245 4.130 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.550 0.995 2.060 ;
        RECT 0.730 0.750 0.995 1.550 ;
        RECT 0.730 0.350 1.060 0.750 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.215 2.570 0.545 3.245 ;
        RECT 1.115 2.570 1.445 3.245 ;
        RECT 1.635 2.570 1.965 2.980 ;
        RECT 2.135 2.740 2.665 3.245 ;
        RECT 2.835 2.570 3.165 2.980 ;
        RECT 0.105 2.230 1.335 2.400 ;
        RECT 1.635 2.290 3.165 2.570 ;
        RECT 0.105 1.350 0.435 2.230 ;
        RECT 1.165 2.120 1.335 2.230 ;
        RECT 3.705 2.120 4.035 2.980 ;
        RECT 1.165 1.950 4.035 2.120 ;
        RECT 0.300 0.085 0.550 1.130 ;
        RECT 1.165 1.090 1.335 1.950 ;
        RECT 1.165 0.920 4.040 1.090 ;
        RECT 1.230 0.085 1.630 0.750 ;
        RECT 2.630 0.350 3.000 0.920 ;
        RECT 3.170 0.085 3.540 0.750 ;
        RECT 3.710 0.350 4.040 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a311o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a311o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a311o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.450 7.075 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 7.245 1.450 7.575 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.420 5.295 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.470 1.865 1.800 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.495 1.470 0.825 1.800 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.275 1.295 7.625 1.355 ;
        RECT 2.990 1.280 7.625 1.295 ;
        RECT 2.085 1.180 7.625 1.280 ;
        RECT 0.305 0.245 7.625 1.180 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER met1 ;
        RECT 0.095 0.995 0.385 1.040 ;
        RECT 2.495 0.995 2.785 1.040 ;
        RECT 0.095 0.855 2.785 0.995 ;
        RECT 0.095 0.810 0.385 0.855 ;
        RECT 2.495 0.810 2.785 0.855 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 1.205 2.980 2.435 3.075 ;
        RECT 0.305 2.905 2.435 2.980 ;
        RECT 0.305 2.700 1.535 2.905 ;
        RECT 0.125 2.360 1.505 2.530 ;
        RECT 0.125 1.040 0.295 2.360 ;
        RECT 0.755 2.020 1.165 2.190 ;
        RECT 0.995 1.300 1.165 2.020 ;
        RECT 1.335 2.140 1.505 2.360 ;
        RECT 1.735 2.490 1.905 2.735 ;
        RECT 2.105 2.660 2.435 2.905 ;
        RECT 2.625 2.660 2.955 3.245 ;
        RECT 3.525 2.660 3.855 3.245 ;
        RECT 4.425 2.660 4.755 3.245 ;
        RECT 4.940 2.490 5.270 2.980 ;
        RECT 5.470 2.630 5.720 3.245 ;
        RECT 1.735 2.460 5.270 2.490 ;
        RECT 5.920 2.460 6.090 2.980 ;
        RECT 1.735 2.320 6.090 2.460 ;
        RECT 1.735 2.310 1.905 2.320 ;
        RECT 4.940 2.290 6.090 2.320 ;
        RECT 6.290 2.290 6.650 3.245 ;
        RECT 2.525 2.140 4.305 2.150 ;
        RECT 1.335 1.970 4.305 2.140 ;
        RECT 5.920 2.120 6.090 2.290 ;
        RECT 6.850 2.120 7.020 2.980 ;
        RECT 2.525 1.820 4.305 1.970 ;
        RECT 4.475 1.950 5.715 2.120 ;
        RECT 5.920 1.950 7.020 2.120 ;
        RECT 7.220 1.950 7.550 3.245 ;
        RECT 4.475 1.650 4.645 1.950 ;
        RECT 2.055 1.480 4.645 1.650 ;
        RECT 2.055 1.320 3.905 1.480 ;
        RECT 2.055 1.300 2.325 1.320 ;
        RECT 0.905 1.130 2.325 1.300 ;
        RECT 5.545 1.265 5.715 1.950 ;
        RECT 4.175 1.150 5.175 1.185 ;
        RECT 0.125 0.810 0.355 1.040 ;
        RECT 0.395 0.085 0.725 0.640 ;
        RECT 0.905 0.390 1.085 1.130 ;
        RECT 1.255 0.085 1.585 0.960 ;
        RECT 1.755 0.390 1.935 1.130 ;
        RECT 2.535 0.980 3.745 1.150 ;
        RECT 2.115 0.085 2.365 0.960 ;
        RECT 2.535 0.390 2.920 0.980 ;
        RECT 3.100 0.085 3.315 0.810 ;
        RECT 3.495 0.405 3.745 0.980 ;
        RECT 3.925 0.935 5.175 1.150 ;
        RECT 5.545 0.935 6.105 1.265 ;
        RECT 6.285 0.985 7.535 1.245 ;
        RECT 3.925 0.085 4.175 0.935 ;
        RECT 6.775 0.765 7.105 0.815 ;
        RECT 4.415 0.595 7.105 0.765 ;
        RECT 4.415 0.505 4.745 0.595 ;
        RECT 7.285 0.425 7.535 0.985 ;
        RECT 5.365 0.255 7.535 0.425 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 0.840 0.325 1.010 ;
        RECT 2.555 0.840 2.725 1.010 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__a311o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a311oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a311oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.350 1.335 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.495 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.755 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.350 3.255 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.250 0.245 3.170 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.792700 ;
    PORT
      LAYER li1 ;
        RECT 2.775 2.120 3.105 2.980 ;
        RECT 0.665 1.950 3.105 2.120 ;
        RECT 0.665 1.180 0.835 1.950 ;
        RECT 0.665 1.010 3.080 1.180 ;
        RECT 1.085 0.350 2.040 1.010 ;
        RECT 2.750 0.350 3.080 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.315 2.290 0.565 3.245 ;
        RECT 0.765 2.460 1.095 2.980 ;
        RECT 1.265 2.630 1.675 3.245 ;
        RECT 1.845 2.460 2.175 2.980 ;
        RECT 0.765 2.290 2.175 2.460 ;
        RECT 0.340 0.085 0.670 0.840 ;
        RECT 2.210 0.085 2.580 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a311oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a311oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a311oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.870 1.550 3.235 1.780 ;
        RECT 2.300 1.350 3.235 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.220 2.090 1.550 ;
        RECT 1.085 1.180 1.315 1.220 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.470 1.220 0.835 1.550 ;
        RECT 0.605 1.180 0.835 1.220 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.675 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 4.845 1.350 5.175 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.095 0.245 5.105 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.935400 ;
    PORT
      LAYER li1 ;
        RECT 4.850 2.120 5.020 2.735 ;
        RECT 4.850 1.950 5.635 2.120 ;
        RECT 5.405 1.180 5.635 1.950 ;
        RECT 2.555 1.010 5.635 1.180 ;
        RECT 2.555 0.850 3.745 1.010 ;
        RECT 3.495 0.350 3.745 0.850 ;
        RECT 4.685 0.350 5.635 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.170 1.820 0.420 3.245 ;
        RECT 0.620 1.890 0.950 2.980 ;
        RECT 1.150 2.060 1.320 3.245 ;
        RECT 1.520 1.890 1.850 2.980 ;
        RECT 2.050 2.060 2.330 3.245 ;
        RECT 2.530 2.120 2.700 2.980 ;
        RECT 2.900 2.290 3.230 3.245 ;
        RECT 3.420 2.905 5.550 3.075 ;
        RECT 3.420 2.290 3.755 2.905 ;
        RECT 3.925 2.120 4.120 2.735 ;
        RECT 2.530 1.950 4.120 2.120 ;
        RECT 4.320 1.950 4.650 2.905 ;
        RECT 5.220 2.290 5.550 2.905 ;
        RECT 2.530 1.890 2.700 1.950 ;
        RECT 0.620 1.720 2.700 1.890 ;
        RECT 0.185 1.010 0.435 1.050 ;
        RECT 1.905 1.010 2.235 1.050 ;
        RECT 0.185 0.840 2.235 1.010 ;
        RECT 0.185 0.350 0.435 0.840 ;
        RECT 1.125 0.770 2.235 0.840 ;
        RECT 0.615 0.085 0.945 0.670 ;
        RECT 1.125 0.330 1.295 0.770 ;
        RECT 2.985 0.600 3.315 0.680 ;
        RECT 1.475 0.350 3.315 0.600 ;
        RECT 3.915 0.085 4.515 0.840 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__a311oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a311oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a311oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.635 1.350 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 3.715 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.350 1.875 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 6.775 1.320 7.785 1.650 ;
        RECT 6.775 1.180 7.555 1.320 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 8.065 1.220 9.075 1.550 ;
        RECT 8.285 1.180 9.075 1.220 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.245 9.060 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.700600 ;
    PORT
      LAYER li1 ;
        RECT 8.355 1.890 8.525 2.735 ;
        RECT 9.255 1.890 9.425 2.735 ;
        RECT 8.355 1.720 9.425 1.890 ;
        RECT 4.330 1.010 6.380 1.130 ;
        RECT 7.760 1.010 8.010 1.050 ;
        RECT 9.255 1.010 9.425 1.720 ;
        RECT 4.330 0.850 9.425 1.010 ;
        RECT 4.330 0.770 4.660 0.850 ;
        RECT 6.130 0.840 9.425 0.850 ;
        RECT 6.130 0.350 6.380 0.840 ;
        RECT 7.760 0.350 8.010 0.840 ;
        RECT 8.700 0.670 9.425 0.840 ;
        RECT 8.700 0.350 9.955 0.670 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.105 1.820 0.355 3.245 ;
        RECT 0.555 2.120 0.805 2.980 ;
        RECT 1.005 2.290 1.335 3.245 ;
        RECT 1.535 2.120 1.705 2.980 ;
        RECT 1.905 2.290 2.235 3.245 ;
        RECT 2.435 2.120 2.605 2.980 ;
        RECT 2.805 2.290 3.135 3.245 ;
        RECT 3.335 2.120 3.505 2.980 ;
        RECT 3.705 2.290 4.035 3.245 ;
        RECT 4.235 2.120 4.405 2.980 ;
        RECT 4.605 2.290 4.855 3.245 ;
        RECT 5.055 2.120 5.305 2.980 ;
        RECT 5.505 2.290 5.835 3.245 ;
        RECT 6.025 2.905 9.955 3.075 ;
        RECT 6.025 2.320 6.355 2.905 ;
        RECT 6.525 2.150 6.755 2.735 ;
        RECT 6.925 2.320 7.255 2.905 ;
        RECT 7.425 2.150 7.655 2.735 ;
        RECT 6.475 2.120 7.655 2.150 ;
        RECT 0.555 1.950 7.655 2.120 ;
        RECT 4.235 1.820 4.405 1.950 ;
        RECT 6.475 1.820 7.655 1.950 ;
        RECT 7.825 1.820 8.155 2.905 ;
        RECT 8.725 2.060 9.055 2.905 ;
        RECT 9.625 1.820 9.955 2.905 ;
        RECT 0.150 1.010 3.920 1.180 ;
        RECT 0.150 0.350 0.400 1.010 ;
        RECT 0.580 0.085 0.830 0.840 ;
        RECT 1.010 0.350 1.260 1.010 ;
        RECT 1.950 0.975 3.920 1.010 ;
        RECT 1.440 0.085 1.770 0.840 ;
        RECT 1.950 0.350 2.120 0.975 ;
        RECT 2.730 0.770 3.060 0.975 ;
        RECT 3.590 0.770 3.920 0.975 ;
        RECT 2.300 0.600 2.560 0.680 ;
        RECT 3.230 0.600 3.420 0.680 ;
        RECT 5.620 0.600 5.950 0.680 ;
        RECT 2.300 0.350 5.950 0.600 ;
        RECT 6.550 0.085 7.590 0.670 ;
        RECT 8.190 0.085 8.520 0.670 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__a311oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a2111o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2111o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.440 0.840 0.670 ;
        RECT 0.510 0.255 0.840 0.440 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.500 2.275 1.800 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.595 0.490 1.795 0.670 ;
        RECT 1.435 0.255 1.795 0.490 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.490 2.245 0.670 ;
        RECT 2.005 0.255 2.335 0.490 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.500 2.775 1.800 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.295 1.260 3.185 1.450 ;
        RECT 0.295 0.245 4.285 1.260 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 3.860 0.370 4.195 2.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.360 2.140 0.690 2.980 ;
        RECT 0.890 2.310 1.100 3.245 ;
        RECT 1.300 2.140 1.630 2.980 ;
        RECT 0.360 1.970 1.630 2.140 ;
        RECT 2.530 2.140 2.860 2.980 ;
        RECT 2.530 1.970 3.115 2.140 ;
        RECT 0.360 1.940 0.690 1.970 ;
        RECT 2.945 1.650 3.115 1.970 ;
        RECT 3.410 1.820 3.660 3.245 ;
        RECT 0.385 1.330 0.715 1.340 ;
        RECT 2.945 1.330 3.690 1.650 ;
        RECT 0.385 1.320 3.690 1.330 ;
        RECT 0.385 1.160 3.115 1.320 ;
        RECT 0.385 0.840 0.715 1.160 ;
        RECT 1.095 0.660 1.425 0.990 ;
        RECT 1.715 0.840 2.045 1.160 ;
        RECT 2.415 0.660 2.675 0.990 ;
        RECT 2.845 0.660 3.115 1.160 ;
        RECT 1.095 0.085 1.265 0.660 ;
        RECT 2.505 0.085 2.675 0.660 ;
        RECT 3.435 0.085 3.685 1.150 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__a2111o_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a2111o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2111o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.350 4.695 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.195 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.350 3.315 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.350 2.775 2.890 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 2.275 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.245 4.610 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.550 0.860 2.980 ;
        RECT 0.690 0.350 0.860 1.550 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.155 1.820 0.405 3.245 ;
        RECT 1.055 2.290 1.385 3.245 ;
        RECT 1.755 2.120 2.085 2.980 ;
        RECT 1.190 1.950 2.085 2.120 ;
        RECT 3.135 2.120 3.505 2.980 ;
        RECT 3.675 2.290 4.045 3.245 ;
        RECT 4.215 2.120 4.545 2.980 ;
        RECT 3.135 1.950 4.545 2.120 ;
        RECT 1.190 1.550 1.360 1.950 ;
        RECT 1.030 1.220 1.360 1.550 ;
        RECT 1.190 1.180 1.360 1.220 ;
        RECT 0.180 0.085 0.510 1.130 ;
        RECT 1.190 1.010 4.520 1.180 ;
        RECT 1.040 0.085 1.370 0.840 ;
        RECT 1.780 0.350 2.030 1.010 ;
        RECT 2.210 0.085 2.580 0.840 ;
        RECT 2.760 0.350 3.010 1.010 ;
        RECT 3.180 0.085 3.730 0.840 ;
        RECT 4.190 0.350 4.520 1.010 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__a2111o_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a2111o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2111o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.285 1.450 7.075 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 7.245 1.260 8.035 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.450 6.115 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.450 5.155 1.780 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.385 1.260 3.715 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.795 1.140 3.030 1.240 ;
        RECT 0.795 0.245 8.150 1.140 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.970 1.165 2.980 ;
        RECT 1.735 1.970 2.065 2.980 ;
        RECT 0.125 1.800 2.065 1.970 ;
        RECT 0.125 1.130 0.650 1.800 ;
        RECT 0.125 0.960 2.445 1.130 ;
        RECT 1.415 0.350 1.665 0.960 ;
        RECT 2.195 0.350 2.445 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.385 2.140 0.635 3.245 ;
        RECT 1.365 2.140 1.535 3.245 ;
        RECT 2.265 1.820 2.515 3.245 ;
        RECT 2.705 2.905 4.835 3.075 ;
        RECT 2.705 2.290 3.035 2.905 ;
        RECT 3.235 2.120 3.405 2.735 ;
        RECT 3.045 1.950 3.405 2.120 ;
        RECT 3.605 1.950 3.935 2.905 ;
        RECT 4.135 2.120 4.305 2.735 ;
        RECT 4.505 2.290 4.835 2.905 ;
        RECT 5.025 2.905 6.175 3.075 ;
        RECT 5.025 2.290 5.305 2.905 ;
        RECT 5.475 2.120 5.805 2.735 ;
        RECT 4.135 1.950 5.805 2.120 ;
        RECT 6.005 2.120 6.175 2.905 ;
        RECT 6.375 2.290 6.705 3.245 ;
        RECT 6.905 2.120 7.075 2.980 ;
        RECT 7.275 2.290 7.525 3.245 ;
        RECT 7.725 2.120 8.055 2.980 ;
        RECT 6.005 1.950 8.055 2.120 ;
        RECT 3.045 1.630 3.215 1.950 ;
        RECT 0.870 1.300 3.215 1.630 ;
        RECT 3.045 1.090 3.215 1.300 ;
        RECT 4.050 1.110 6.770 1.280 ;
        RECT 4.050 1.090 4.220 1.110 ;
        RECT 0.905 0.085 1.235 0.790 ;
        RECT 1.845 0.085 2.015 0.790 ;
        RECT 2.625 0.085 2.875 1.030 ;
        RECT 3.045 0.920 4.220 1.090 ;
        RECT 3.045 0.350 3.350 0.920 ;
        RECT 3.530 0.085 3.870 0.750 ;
        RECT 4.050 0.350 4.220 0.920 ;
        RECT 4.400 0.085 4.740 0.940 ;
        RECT 4.920 0.350 5.090 1.110 ;
        RECT 5.270 0.085 5.600 0.940 ;
        RECT 6.010 0.455 6.340 0.940 ;
        RECT 6.510 0.625 6.770 1.110 ;
        RECT 6.950 0.920 8.060 1.090 ;
        RECT 6.950 0.455 7.120 0.920 ;
        RECT 6.010 0.285 7.120 0.455 ;
        RECT 7.300 0.085 7.630 0.750 ;
        RECT 7.810 0.350 8.060 0.920 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__a2111o_4

#--------EOF---------

MACRO sky130_fd_sc_hs__a2111oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2111oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.415 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.625 1.180 3.235 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.350 1.335 1.780 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.465 1.350 0.835 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.250 0.245 3.190 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.950 1.315 2.980 ;
        RECT 0.125 1.180 0.295 1.950 ;
        RECT 0.125 1.010 2.180 1.180 ;
        RECT 0.850 0.350 1.100 1.010 ;
        RECT 1.850 0.350 2.180 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 1.695 2.120 2.065 2.980 ;
        RECT 2.235 2.290 2.605 3.245 ;
        RECT 2.775 2.120 3.105 2.980 ;
        RECT 1.695 1.950 3.105 2.120 ;
        RECT 2.775 1.820 3.105 1.950 ;
        RECT 0.340 0.085 0.670 0.840 ;
        RECT 1.270 0.085 1.680 0.840 ;
        RECT 2.750 0.085 3.080 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__a2111oi_1

#--------EOF---------

MACRO sky130_fd_sc_hs__a2111oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2111oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 4.675 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.850 1.350 5.180 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.180 3.715 1.550 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.350 2.755 1.780 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 1.315 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.550 0.245 2.590 1.240 ;
        RECT 3.480 0.245 5.720 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.027900 ;
    PORT
      LAYER li1 ;
        RECT 0.755 2.120 1.085 2.735 ;
        RECT 0.125 1.950 1.085 2.120 ;
        RECT 0.125 1.180 0.355 1.950 ;
        RECT 0.125 1.010 2.500 1.180 ;
        RECT 1.160 0.350 1.490 1.010 ;
        RECT 2.170 0.975 2.500 1.010 ;
        RECT 4.000 0.975 4.330 1.130 ;
        RECT 2.170 0.770 4.330 0.975 ;
        RECT 2.170 0.350 2.500 0.770 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.305 2.905 2.435 3.075 ;
        RECT 0.305 2.290 0.555 2.905 ;
        RECT 1.285 1.950 1.455 2.905 ;
        RECT 1.655 2.120 1.985 2.735 ;
        RECT 2.185 2.290 2.435 2.905 ;
        RECT 2.625 2.905 3.855 3.075 ;
        RECT 2.625 2.290 2.905 2.905 ;
        RECT 3.075 2.120 3.325 2.735 ;
        RECT 1.655 1.950 3.325 2.120 ;
        RECT 3.525 2.120 3.855 2.905 ;
        RECT 4.055 2.290 4.225 3.245 ;
        RECT 4.425 2.120 4.675 2.980 ;
        RECT 4.875 2.290 5.205 3.245 ;
        RECT 5.405 2.120 5.655 2.980 ;
        RECT 3.525 1.950 5.655 2.120 ;
        RECT 3.075 1.820 3.325 1.950 ;
        RECT 5.405 1.820 5.655 1.950 ;
        RECT 4.510 1.010 5.630 1.180 ;
        RECT 0.660 0.085 0.990 0.840 ;
        RECT 1.660 0.085 2.000 0.840 ;
        RECT 4.510 0.600 4.680 1.010 ;
        RECT 3.570 0.350 4.680 0.600 ;
        RECT 4.860 0.085 5.200 0.840 ;
        RECT 5.380 0.350 5.630 1.010 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__a2111oi_2

#--------EOF---------

MACRO sky130_fd_sc_hs__a2111oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a2111oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.450 1.350 8.035 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.205 1.350 9.555 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.350 6.075 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 2.235 1.350 3.510 1.780 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.180 1.905 1.550 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.930 0.245 4.920 1.240 ;
        RECT 6.010 0.245 10.000 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.708000 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.890 0.885 2.735 ;
        RECT 1.455 1.890 1.705 2.735 ;
        RECT 0.125 1.720 1.705 1.890 ;
        RECT 0.125 1.010 0.355 1.720 ;
        RECT 2.390 1.130 6.880 1.180 ;
        RECT 2.390 1.010 7.740 1.130 ;
        RECT 0.125 0.840 2.640 1.010 ;
        RECT 1.530 0.330 1.700 0.840 ;
        RECT 2.390 0.350 2.640 0.840 ;
        RECT 4.070 0.975 7.740 1.010 ;
        RECT 4.070 0.350 4.320 0.975 ;
        RECT 6.550 0.915 7.740 0.975 ;
        RECT 6.550 0.770 6.880 0.915 ;
        RECT 7.410 0.770 7.740 0.915 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.105 2.905 2.235 3.075 ;
        RECT 0.105 2.060 0.355 2.905 ;
        RECT 1.085 2.060 1.255 2.905 ;
        RECT 1.905 2.120 2.235 2.905 ;
        RECT 2.435 2.905 5.925 3.075 ;
        RECT 2.435 2.290 2.685 2.905 ;
        RECT 2.855 2.120 3.085 2.735 ;
        RECT 3.255 2.290 3.585 2.905 ;
        RECT 3.755 2.120 4.035 2.735 ;
        RECT 1.905 1.950 4.035 2.120 ;
        RECT 4.245 2.120 4.525 2.735 ;
        RECT 4.695 2.290 5.025 2.905 ;
        RECT 5.195 2.120 5.425 2.735 ;
        RECT 5.595 2.290 5.925 2.905 ;
        RECT 6.125 2.120 6.295 2.980 ;
        RECT 6.495 2.290 6.825 3.245 ;
        RECT 7.025 2.120 7.195 2.980 ;
        RECT 7.395 2.290 7.725 3.245 ;
        RECT 7.925 2.120 8.095 2.980 ;
        RECT 8.295 2.290 8.545 3.245 ;
        RECT 8.745 2.120 9.075 2.980 ;
        RECT 9.275 2.290 9.525 3.245 ;
        RECT 9.725 2.120 9.975 2.980 ;
        RECT 4.245 1.950 9.975 2.120 ;
        RECT 3.705 1.820 4.035 1.950 ;
        RECT 9.725 1.820 9.975 1.950 ;
        RECT 7.920 1.010 9.890 1.180 ;
        RECT 1.020 0.085 1.350 0.670 ;
        RECT 1.880 0.085 2.210 0.670 ;
        RECT 2.810 0.085 3.900 0.840 ;
        RECT 4.500 0.085 4.830 0.805 ;
        RECT 6.120 0.600 6.380 0.680 ;
        RECT 7.040 0.600 7.250 0.680 ;
        RECT 7.920 0.600 8.090 1.010 ;
        RECT 6.120 0.350 8.090 0.600 ;
        RECT 8.270 0.085 8.600 0.840 ;
        RECT 8.780 0.350 8.950 1.010 ;
        RECT 9.130 0.085 9.460 0.840 ;
        RECT 9.640 0.350 9.890 1.010 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__a2111oi_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 0.835 0.670 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.075 1.180 1.405 1.680 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 1.370 1.095 1.450 ;
        RECT 0.150 0.245 2.280 1.370 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 1.920 1.850 2.315 2.980 ;
        RECT 2.145 1.180 2.315 1.850 ;
        RECT 1.840 0.470 2.315 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.350 2.190 0.685 3.245 ;
        RECT 0.855 2.020 1.185 3.000 ;
        RECT 1.390 2.190 1.720 3.245 ;
        RECT 0.260 1.850 1.750 2.020 ;
        RECT 0.260 0.840 0.590 1.850 ;
        RECT 1.580 1.680 1.750 1.850 ;
        RECT 1.580 1.350 1.975 1.680 ;
        RECT 1.340 0.085 1.670 1.010 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__and2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.300 1.085 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.595 1.890 1.845 2.980 ;
        RECT 1.595 1.720 2.010 1.890 ;
        RECT 1.840 1.020 2.010 1.720 ;
        RECT 1.625 0.850 2.010 1.020 ;
        RECT 1.625 0.790 1.795 0.850 ;
        RECT 1.465 0.350 1.795 0.790 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.110 1.950 0.440 3.245 ;
        RECT 0.640 2.120 0.890 2.980 ;
        RECT 1.060 2.290 1.390 3.245 ;
        RECT 0.640 1.950 1.425 2.120 ;
        RECT 2.045 2.060 2.295 3.245 ;
        RECT 1.255 1.550 1.425 1.950 ;
        RECT 1.255 1.220 1.670 1.550 ;
        RECT 1.255 1.130 1.425 1.220 ;
        RECT 0.135 0.960 1.425 1.130 ;
        RECT 0.135 0.350 0.465 0.960 ;
        RECT 0.955 0.085 1.285 0.790 ;
        RECT 1.975 0.085 2.285 0.680 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__and2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.450 3.255 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 2.255 1.345 2.755 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.315 1.365 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.219800 ;
    PORT
      LAYER li1 ;
        RECT 0.545 2.015 0.815 2.980 ;
        RECT 1.465 2.015 1.715 2.980 ;
        RECT 0.545 1.845 1.715 2.015 ;
        RECT 0.545 1.550 0.835 1.845 ;
        RECT 0.545 1.175 0.795 1.550 ;
        RECT 0.545 1.005 1.725 1.175 ;
        RECT 0.545 0.475 0.795 1.005 ;
        RECT 1.475 0.475 1.725 1.005 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.015 2.185 1.265 3.245 ;
        RECT 1.935 2.290 2.265 3.245 ;
        RECT 2.470 2.120 2.800 2.905 ;
        RECT 2.970 2.290 3.300 3.245 ;
        RECT 3.500 2.120 3.670 2.905 ;
        RECT 1.885 1.950 3.670 2.120 ;
        RECT 3.870 2.025 4.200 3.245 ;
        RECT 1.885 1.675 2.055 1.950 ;
        RECT 1.005 1.345 2.055 1.675 ;
        RECT 3.500 1.280 3.670 1.950 ;
        RECT 0.115 0.085 0.365 1.255 ;
        RECT 0.975 0.085 1.305 0.835 ;
        RECT 1.985 0.085 2.315 1.175 ;
        RECT 2.495 0.425 2.825 1.175 ;
        RECT 2.995 1.110 3.670 1.280 ;
        RECT 2.995 0.595 3.325 1.110 ;
        RECT 3.505 0.425 3.675 0.940 ;
        RECT 2.495 0.255 3.675 0.425 ;
        RECT 3.875 0.085 4.205 1.255 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__and2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 2.150 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.375 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.200 1.050 3.355 1.260 ;
        RECT 0.005 0.245 3.355 1.050 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 2.770 1.820 3.255 2.980 ;
        RECT 3.085 1.150 3.255 1.820 ;
        RECT 2.915 0.370 3.255 1.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.320 1.165 2.650 ;
        RECT 0.810 1.180 1.140 2.320 ;
        RECT 1.365 1.820 1.535 3.245 ;
        RECT 1.705 1.950 2.065 2.700 ;
        RECT 2.270 1.950 2.600 3.245 ;
        RECT 0.115 1.010 1.140 1.180 ;
        RECT 1.705 1.150 1.875 1.950 ;
        RECT 2.575 1.320 2.915 1.650 ;
        RECT 2.575 1.150 2.745 1.320 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 1.310 0.980 2.745 1.150 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.310 0.470 1.640 0.980 ;
        RECT 2.130 0.085 2.745 0.810 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__and2b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.525 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.610 1.050 3.330 1.240 ;
        RECT 0.005 0.245 3.330 1.050 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.820 1.515 2.150 ;
        RECT 1.115 1.130 1.285 1.820 ;
        RECT 1.115 0.350 1.445 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.490 0.445 2.700 ;
        RECT 0.650 2.660 0.980 3.245 ;
        RECT 1.635 2.660 2.260 3.245 ;
        RECT 2.915 2.660 3.245 3.245 ;
        RECT 0.115 2.320 3.135 2.490 ;
        RECT 0.115 1.950 0.890 2.320 ;
        RECT 0.720 1.180 0.890 1.950 ;
        RECT 1.685 1.870 2.795 2.150 ;
        RECT 1.685 1.630 1.855 1.870 ;
        RECT 2.965 1.630 3.135 2.320 ;
        RECT 1.455 1.300 1.855 1.630 ;
        RECT 2.765 1.300 3.135 1.630 ;
        RECT 0.115 1.010 0.890 1.180 ;
        RECT 1.685 1.010 1.855 1.300 ;
        RECT 2.890 1.010 3.220 1.130 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 1.685 0.840 3.220 1.010 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.615 0.085 2.400 0.600 ;
        RECT 2.890 0.350 3.220 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__and2b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.450 0.805 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.620 2.585 1.790 ;
        RECT 0.975 1.435 1.305 1.620 ;
        RECT 2.045 1.180 2.585 1.620 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.500 1.140 4.780 1.240 ;
        RECT 0.100 0.245 4.780 1.140 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.093800 ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.990 3.265 2.980 ;
        RECT 3.995 1.990 4.165 2.980 ;
        RECT 3.095 1.820 4.165 1.990 ;
        RECT 3.995 1.650 4.165 1.820 ;
        RECT 3.995 1.480 4.675 1.650 ;
        RECT 4.445 1.150 4.675 1.480 ;
        RECT 3.095 0.980 4.675 1.150 ;
        RECT 3.095 0.350 3.265 0.980 ;
        RECT 3.910 0.350 4.160 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.085 1.950 0.355 2.980 ;
        RECT 0.555 2.100 0.885 3.245 ;
        RECT 1.075 2.130 1.405 2.980 ;
        RECT 1.605 2.300 1.855 3.245 ;
        RECT 2.045 2.130 2.375 2.980 ;
        RECT 2.565 2.300 2.895 3.245 ;
        RECT 3.465 2.160 3.795 3.245 ;
        RECT 1.075 1.960 2.925 2.130 ;
        RECT 0.085 1.265 0.255 1.950 ;
        RECT 2.755 1.650 2.925 1.960 ;
        RECT 4.365 1.820 4.695 3.245 ;
        RECT 1.515 1.265 1.845 1.450 ;
        RECT 0.085 1.095 1.845 1.265 ;
        RECT 2.755 1.320 3.825 1.650 ;
        RECT 0.085 0.350 0.540 1.095 ;
        RECT 2.755 0.925 2.925 1.320 ;
        RECT 0.710 0.085 1.040 0.925 ;
        RECT 1.210 0.585 1.470 0.925 ;
        RECT 1.640 0.755 2.925 0.925 ;
        RECT 1.210 0.335 2.400 0.585 ;
        RECT 2.570 0.085 2.900 0.585 ;
        RECT 3.445 0.085 3.695 0.810 ;
        RECT 4.340 0.085 4.670 0.810 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__and2b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.570 1.315 0.670 ;
        RECT 0.105 0.255 1.315 0.570 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.180 1.315 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.450 1.815 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 1.370 1.545 1.450 ;
        RECT 0.040 0.245 2.635 1.370 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 2.480 1.850 2.765 2.980 ;
        RECT 2.595 1.180 2.765 1.850 ;
        RECT 2.195 1.010 2.765 1.180 ;
        RECT 2.195 0.480 2.525 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.115 2.120 0.445 2.850 ;
        RECT 0.615 2.290 0.945 3.245 ;
        RECT 1.115 2.120 1.400 2.850 ;
        RECT 1.570 2.290 2.310 3.245 ;
        RECT 0.115 1.950 2.240 2.120 ;
        RECT 0.115 0.740 0.480 1.950 ;
        RECT 2.070 1.680 2.240 1.950 ;
        RECT 2.070 1.350 2.400 1.680 ;
        RECT 1.695 0.085 2.025 1.180 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__and3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.255 1.315 0.670 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.905 1.180 1.315 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.430 1.815 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 1.280 2.005 1.450 ;
        RECT 0.100 0.245 3.285 1.280 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.572800 ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.840 2.725 2.980 ;
        RECT 2.555 1.170 2.725 1.840 ;
        RECT 2.180 0.810 2.755 1.170 ;
        RECT 2.180 0.390 2.510 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.185 2.120 0.515 2.780 ;
        RECT 0.685 2.290 1.015 3.245 ;
        RECT 1.205 2.120 1.535 2.780 ;
        RECT 1.875 2.290 2.205 3.245 ;
        RECT 0.185 1.950 2.205 2.120 ;
        RECT 0.185 1.340 0.515 1.950 ;
        RECT 2.035 1.670 2.205 1.950 ;
        RECT 2.895 1.820 3.225 3.245 ;
        RECT 2.035 1.340 2.385 1.670 ;
        RECT 0.185 0.840 0.540 1.340 ;
        RECT 1.680 0.085 2.010 1.170 ;
        RECT 2.925 0.640 3.245 1.170 ;
        RECT 2.680 0.085 3.245 0.640 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__and3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 4.615 1.450 5.285 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.325 4.335 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.450 3.230 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 1.140 2.325 1.240 ;
        RECT 0.020 0.245 5.750 1.140 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.970 0.895 2.980 ;
        RECT 1.565 1.970 1.895 2.980 ;
        RECT 0.560 1.800 1.895 1.970 ;
        RECT 0.560 1.130 0.835 1.800 ;
        RECT 0.560 0.960 1.740 1.130 ;
        RECT 0.560 0.350 0.890 0.960 ;
        RECT 1.490 0.350 1.740 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.065 2.140 1.395 3.245 ;
        RECT 2.065 2.290 2.395 3.245 ;
        RECT 2.565 2.120 2.895 2.980 ;
        RECT 3.065 2.290 3.645 3.245 ;
        RECT 3.815 2.120 4.145 2.980 ;
        RECT 4.315 2.290 4.645 3.245 ;
        RECT 4.815 2.120 5.145 2.980 ;
        RECT 5.315 2.290 5.645 3.245 ;
        RECT 2.065 1.950 5.625 2.120 ;
        RECT 2.065 1.630 2.235 1.950 ;
        RECT 1.035 1.300 2.235 1.630 ;
        RECT 5.455 1.280 5.625 1.950 ;
        RECT 0.130 0.085 0.380 1.130 ;
        RECT 1.070 0.085 1.320 0.790 ;
        RECT 1.920 0.085 2.250 1.030 ;
        RECT 2.420 0.985 4.090 1.155 ;
        RECT 4.810 1.110 5.625 1.280 ;
        RECT 2.420 0.350 2.670 0.985 ;
        RECT 2.850 0.085 3.180 0.815 ;
        RECT 3.410 0.425 3.740 0.815 ;
        RECT 3.920 0.595 4.090 0.985 ;
        RECT 4.310 0.425 4.640 1.030 ;
        RECT 4.810 0.595 5.140 1.110 ;
        RECT 5.310 0.425 5.640 0.940 ;
        RECT 3.410 0.255 5.640 0.425 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__and3_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.110 0.570 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.005 1.390 2.335 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.390 2.875 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.200 1.050 3.825 1.240 ;
        RECT 0.005 0.245 3.825 1.050 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.345 1.820 3.755 2.980 ;
        RECT 3.585 1.130 3.755 1.820 ;
        RECT 3.385 0.350 3.755 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 2.100 0.445 3.245 ;
        RECT 0.615 2.100 0.945 2.980 ;
        RECT 0.775 1.700 0.945 2.100 ;
        RECT 1.310 2.120 1.640 2.700 ;
        RECT 1.810 2.290 2.140 3.245 ;
        RECT 2.310 2.120 2.640 2.700 ;
        RECT 1.310 1.950 2.640 2.120 ;
        RECT 2.845 1.950 3.175 3.245 ;
        RECT 0.775 1.030 1.140 1.700 ;
        RECT 1.310 1.220 1.640 1.950 ;
        RECT 3.045 1.300 3.415 1.630 ;
        RECT 3.045 1.220 3.215 1.300 ;
        RECT 1.310 1.050 3.215 1.220 ;
        RECT 0.775 0.940 0.945 1.030 ;
        RECT 0.115 0.085 0.445 0.940 ;
        RECT 0.615 0.350 0.945 0.940 ;
        RECT 1.310 0.450 1.640 1.050 ;
        RECT 2.625 0.085 3.215 0.880 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__and3b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.260 0.550 1.930 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.440 2.450 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.690 1.350 3.235 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.315 1.120 4.255 1.240 ;
        RECT 0.005 0.245 4.255 1.120 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.560000 ;
    PORT
      LAYER li1 ;
        RECT 3.410 1.820 3.755 2.070 ;
        RECT 3.410 1.130 3.715 1.820 ;
        RECT 3.385 0.350 3.715 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.270 0.400 2.980 ;
        RECT 0.570 2.440 0.900 3.245 ;
        RECT 0.115 2.100 1.070 2.270 ;
        RECT 0.900 1.855 1.070 2.100 ;
        RECT 1.400 2.120 1.730 2.860 ;
        RECT 1.900 2.290 2.230 3.245 ;
        RECT 2.420 2.410 2.750 2.860 ;
        RECT 2.960 2.580 3.290 3.245 ;
        RECT 3.875 2.580 4.205 3.245 ;
        RECT 2.420 2.240 4.215 2.410 ;
        RECT 2.420 2.120 2.750 2.240 ;
        RECT 1.400 1.950 2.750 2.120 ;
        RECT 0.900 1.090 1.230 1.855 ;
        RECT 0.115 0.920 1.230 1.090 ;
        RECT 0.115 0.420 0.375 0.920 ;
        RECT 0.545 0.085 0.875 0.750 ;
        RECT 1.400 0.350 1.755 1.950 ;
        RECT 4.045 1.630 4.215 2.240 ;
        RECT 3.885 1.300 4.215 1.630 ;
        RECT 2.815 0.085 3.145 1.130 ;
        RECT 3.895 0.085 4.145 1.130 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__and3b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.180 0.835 1.510 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.755 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 3.560 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065 1.240 3.405 1.260 ;
        RECT 1.065 1.140 6.715 1.240 ;
        RECT 0.005 0.245 6.715 1.140 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.138200 ;
    PORT
      LAYER li1 ;
        RECT 4.570 1.970 4.900 2.980 ;
        RECT 5.570 1.970 5.900 2.980 ;
        RECT 4.570 1.800 6.595 1.970 ;
        RECT 5.935 1.130 6.105 1.800 ;
        RECT 6.365 1.550 6.595 1.800 ;
        RECT 4.965 0.960 6.105 1.130 ;
        RECT 4.965 0.350 5.215 0.960 ;
        RECT 5.925 0.350 6.105 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.475 1.850 0.805 2.860 ;
        RECT 0.975 2.020 1.305 3.245 ;
        RECT 1.475 2.120 1.805 2.860 ;
        RECT 1.975 2.290 2.305 3.245 ;
        RECT 2.475 2.120 2.805 2.860 ;
        RECT 2.975 2.290 3.305 3.245 ;
        RECT 3.535 2.120 3.900 2.860 ;
        RECT 1.475 1.950 3.900 2.120 ;
        RECT 0.115 1.680 1.305 1.850 ;
        RECT 1.475 1.820 1.865 1.950 ;
        RECT 0.115 1.010 0.285 1.680 ;
        RECT 1.135 1.650 1.305 1.680 ;
        RECT 1.135 1.320 1.525 1.650 ;
        RECT 1.695 1.150 1.865 1.820 ;
        RECT 3.730 1.630 3.900 1.950 ;
        RECT 4.070 1.820 4.400 3.245 ;
        RECT 5.070 2.140 5.400 3.245 ;
        RECT 6.070 2.140 6.400 3.245 ;
        RECT 3.730 1.460 5.765 1.630 ;
        RECT 4.755 1.300 5.765 1.460 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.875 1.010 ;
        RECT 1.175 0.425 1.505 1.150 ;
        RECT 1.685 0.595 1.865 1.150 ;
        RECT 2.035 0.720 2.365 1.150 ;
        RECT 2.535 1.010 4.285 1.180 ;
        RECT 2.535 0.890 2.865 1.010 ;
        RECT 2.035 0.470 3.295 0.720 ;
        RECT 2.035 0.425 2.365 0.470 ;
        RECT 1.175 0.255 2.365 0.425 ;
        RECT 3.525 0.085 3.855 0.840 ;
        RECT 4.035 0.450 4.285 1.010 ;
        RECT 4.465 0.085 4.795 1.130 ;
        RECT 5.395 0.085 5.725 0.790 ;
        RECT 6.275 0.085 6.605 1.130 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__and3b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.120 0.815 1.790 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.440 1.315 1.805 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.440 1.855 1.790 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.395 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.225 1.140 3.170 1.240 ;
        RECT 0.350 0.245 3.170 1.140 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 2.910 1.820 3.275 2.980 ;
        RECT 3.105 1.130 3.275 1.820 ;
        RECT 2.730 0.350 3.275 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.315 0.445 3.245 ;
        RECT 0.615 2.145 0.945 2.980 ;
        RECT 1.115 2.315 1.705 3.245 ;
        RECT 1.875 2.145 2.205 2.980 ;
        RECT 2.410 2.300 2.740 3.245 ;
        RECT 0.085 2.130 2.205 2.145 ;
        RECT 0.085 1.975 2.740 2.130 ;
        RECT 0.085 0.950 0.255 1.975 ;
        RECT 1.875 1.960 2.740 1.975 ;
        RECT 2.570 1.650 2.740 1.960 ;
        RECT 2.570 1.320 2.935 1.650 ;
        RECT 0.085 0.355 0.770 0.950 ;
        RECT 2.220 0.085 2.550 1.030 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__and4_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.300 0.445 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.440 1.315 1.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.440 1.855 1.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.425 1.550 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 0.245 3.745 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.130 3.235 2.150 ;
        RECT 2.790 0.770 3.235 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 1.950 0.445 3.245 ;
        RECT 0.615 1.890 0.985 2.980 ;
        RECT 1.215 2.060 1.545 3.245 ;
        RECT 1.765 2.490 2.095 2.980 ;
        RECT 2.300 2.660 2.630 3.245 ;
        RECT 3.370 2.660 3.725 3.245 ;
        RECT 1.765 2.320 3.735 2.490 ;
        RECT 1.765 1.890 2.095 2.320 ;
        RECT 0.615 1.720 2.095 1.890 ;
        RECT 0.615 1.130 0.785 1.720 ;
        RECT 3.405 1.300 3.735 2.320 ;
        RECT 0.260 0.960 0.785 1.130 ;
        RECT 0.260 0.350 0.590 0.960 ;
        RECT 2.265 0.085 2.595 1.010 ;
        RECT 3.405 0.600 3.655 1.080 ;
        RECT 3.220 0.085 3.655 0.600 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__and4_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.450 1.390 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.550 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.980 1.345 4.365 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.930 1.470 3.260 1.800 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 1.240 4.180 1.365 ;
        RECT 0.030 0.245 6.635 1.240 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.164600 ;
    PORT
      LAYER li1 ;
        RECT 4.875 1.970 5.205 2.980 ;
        RECT 5.855 1.970 6.105 2.980 ;
        RECT 4.875 1.800 6.105 1.970 ;
        RECT 5.855 1.650 6.105 1.800 ;
        RECT 5.855 1.480 6.595 1.650 ;
        RECT 6.365 1.130 6.595 1.480 ;
        RECT 4.830 0.960 6.595 1.130 ;
        RECT 4.830 0.350 5.080 0.960 ;
        RECT 5.760 0.350 6.090 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.115 1.950 0.395 3.245 ;
        RECT 1.015 2.410 1.345 3.245 ;
        RECT 1.560 2.240 1.730 2.980 ;
        RECT 0.565 1.950 1.730 2.240 ;
        RECT 0.720 1.255 0.890 1.950 ;
        RECT 1.560 1.770 1.730 1.950 ;
        RECT 1.930 1.940 2.260 3.245 ;
        RECT 2.430 2.140 2.760 2.980 ;
        RECT 2.930 2.310 3.645 3.245 ;
        RECT 3.815 2.140 4.145 2.980 ;
        RECT 4.315 2.290 4.645 3.245 ;
        RECT 5.405 2.140 5.655 3.245 ;
        RECT 2.430 2.120 4.145 2.140 ;
        RECT 2.430 1.970 4.705 2.120 ;
        RECT 2.430 1.770 2.760 1.970 ;
        RECT 3.815 1.950 4.705 1.970 ;
        RECT 1.560 1.600 2.760 1.770 ;
        RECT 4.535 1.630 4.705 1.950 ;
        RECT 6.275 1.820 6.605 3.245 ;
        RECT 4.535 1.300 5.685 1.630 ;
        RECT 0.140 0.485 0.390 1.255 ;
        RECT 0.720 1.005 1.330 1.255 ;
        RECT 1.940 1.175 3.810 1.300 ;
        RECT 1.940 1.130 4.070 1.175 ;
        RECT 0.570 0.655 1.760 0.835 ;
        RECT 1.940 0.485 2.110 1.130 ;
        RECT 3.640 0.995 4.070 1.130 ;
        RECT 2.290 0.825 3.470 0.960 ;
        RECT 2.290 0.790 3.640 0.825 ;
        RECT 2.290 0.575 2.620 0.790 ;
        RECT 0.140 0.315 2.110 0.485 ;
        RECT 2.800 0.085 3.130 0.620 ;
        RECT 3.300 0.575 3.640 0.790 ;
        RECT 4.330 0.085 4.660 1.130 ;
        RECT 5.260 0.085 5.590 0.790 ;
        RECT 6.260 0.085 6.520 0.680 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__and4_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.190 0.595 1.860 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.550 2.275 1.960 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.255 2.810 0.670 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.550 3.315 1.880 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.710 1.390 3.010 1.465 ;
        RECT 1.200 1.370 3.010 1.390 ;
        RECT 1.200 1.050 4.315 1.370 ;
        RECT 0.005 0.245 4.315 1.050 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.940 4.510 3.520 ;
        RECT -0.190 1.660 1.370 1.940 ;
        RECT 3.220 1.660 4.510 1.940 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.875 1.850 4.230 2.980 ;
        RECT 4.060 1.180 4.230 1.850 ;
        RECT 3.875 0.480 4.230 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.200 0.445 2.980 ;
        RECT 0.615 2.370 0.945 3.245 ;
        RECT 1.645 2.535 2.595 3.245 ;
        RECT 1.115 2.350 1.460 2.460 ;
        RECT 2.765 2.350 3.095 2.980 ;
        RECT 0.115 2.030 0.945 2.200 ;
        RECT 1.115 2.130 3.095 2.350 ;
        RECT 0.775 1.880 0.945 2.030 ;
        RECT 2.595 2.100 3.095 2.130 ;
        RECT 3.335 2.100 3.665 3.245 ;
        RECT 0.775 1.550 1.255 1.880 ;
        RECT 0.775 1.020 0.945 1.550 ;
        RECT 2.595 1.380 2.765 2.100 ;
        RECT 3.535 1.380 3.890 1.680 ;
        RECT 0.115 0.850 0.945 1.020 ;
        RECT 1.310 1.350 3.890 1.380 ;
        RECT 1.310 1.210 3.705 1.350 ;
        RECT 0.115 0.350 0.405 0.850 ;
        RECT 0.575 0.085 0.875 0.680 ;
        RECT 1.310 0.600 1.640 1.210 ;
        RECT 3.375 0.085 3.705 1.040 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__and4b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 3.405 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.350 2.835 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.350 2.295 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.180 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.820 1.440 2.200 ;
        RECT 1.055 1.130 1.225 1.820 ;
        RECT 1.055 0.350 1.385 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.650 2.710 0.980 3.245 ;
        RECT 1.645 2.710 1.975 3.245 ;
        RECT 2.740 2.710 3.070 3.245 ;
        RECT 3.850 2.710 4.205 3.245 ;
        RECT 0.115 2.540 0.445 2.700 ;
        RECT 0.115 2.370 3.985 2.540 ;
        RECT 0.115 1.950 0.795 2.370 ;
        RECT 0.625 1.130 0.795 1.950 ;
        RECT 1.610 1.950 3.645 2.200 ;
        RECT 1.610 1.630 1.780 1.950 ;
        RECT 3.815 1.680 3.985 2.370 ;
        RECT 1.395 1.300 1.780 1.630 ;
        RECT 3.615 1.350 3.985 1.680 ;
        RECT 0.115 0.960 0.795 1.130 ;
        RECT 1.610 1.130 1.780 1.300 ;
        RECT 1.610 0.960 4.070 1.130 ;
        RECT 0.115 0.540 0.445 0.960 ;
        RECT 0.625 0.085 0.875 0.790 ;
        RECT 1.555 0.085 2.165 0.790 ;
        RECT 3.740 0.350 4.070 0.960 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__and4b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.190 0.835 1.550 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.470 7.180 1.800 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.915 1.350 3.245 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.470 5.155 1.800 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.225 1.290 7.600 1.395 ;
        RECT 3.190 1.240 7.600 1.290 ;
        RECT 0.045 0.245 7.600 1.240 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.209600 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.820 2.405 2.220 ;
        RECT 1.085 1.150 1.315 1.820 ;
        RECT 1.085 0.980 2.540 1.150 ;
        RECT 1.085 0.350 1.470 0.980 ;
        RECT 2.210 0.350 2.540 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.085 2.560 0.445 2.860 ;
        RECT 0.650 2.730 1.025 3.245 ;
        RECT 1.595 2.730 1.955 3.245 ;
        RECT 2.635 2.730 2.980 3.245 ;
        RECT 3.720 2.730 4.050 3.245 ;
        RECT 5.180 2.730 5.530 3.245 ;
        RECT 6.100 2.730 6.430 3.245 ;
        RECT 7.000 2.730 7.565 3.245 ;
        RECT 0.085 2.390 7.520 2.560 ;
        RECT 0.085 1.820 0.445 2.390 ;
        RECT 2.575 1.970 6.880 2.220 ;
        RECT 2.575 1.950 3.515 1.970 ;
        RECT 0.085 1.020 0.255 1.820 ;
        RECT 2.575 1.650 2.745 1.950 ;
        RECT 5.650 1.940 6.080 1.970 ;
        RECT 1.485 1.320 2.745 1.650 ;
        RECT 5.910 1.300 6.080 1.940 ;
        RECT 6.250 1.470 6.675 1.800 ;
        RECT 6.505 1.300 6.675 1.470 ;
        RECT 7.350 1.300 7.520 2.390 ;
        RECT 3.460 1.180 5.475 1.300 ;
        RECT 3.300 1.130 5.475 1.180 ;
        RECT 5.910 1.130 6.335 1.300 ;
        RECT 6.505 1.130 7.520 1.300 ;
        RECT 0.085 0.450 0.405 1.020 ;
        RECT 0.585 0.085 0.915 1.020 ;
        RECT 1.670 0.085 2.000 0.810 ;
        RECT 2.710 0.085 3.040 1.130 ;
        RECT 3.300 0.605 3.630 1.130 ;
        RECT 3.810 0.790 5.125 0.960 ;
        RECT 3.810 0.630 4.105 0.790 ;
        RECT 4.285 0.085 4.615 0.620 ;
        RECT 4.795 0.605 5.125 0.790 ;
        RECT 5.305 0.425 5.475 1.130 ;
        RECT 5.655 0.765 5.905 0.960 ;
        RECT 6.080 0.935 6.335 1.130 ;
        RECT 6.625 0.765 6.955 0.935 ;
        RECT 5.655 0.595 6.955 0.765 ;
        RECT 7.165 0.425 7.495 0.960 ;
        RECT 5.305 0.255 7.495 0.425 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__and4b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.400 1.780 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 4.400 1.300 4.695 1.780 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 3.015 1.190 3.345 1.860 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.190 3.890 1.860 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.515 1.140 1.460 1.240 ;
        RECT 0.515 1.050 4.795 1.140 ;
        RECT 0.005 0.245 4.795 1.050 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.692500 ;
    PORT
      LAYER li1 ;
        RECT 0.910 1.820 1.565 2.150 ;
        RECT 0.910 1.130 1.080 1.820 ;
        RECT 0.910 0.960 1.270 1.130 ;
        RECT 1.080 0.350 1.270 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 2.490 0.445 2.700 ;
        RECT 0.650 2.660 0.980 3.245 ;
        RECT 1.795 2.660 2.125 3.245 ;
        RECT 0.115 2.320 2.045 2.490 ;
        RECT 0.115 1.950 0.740 2.320 ;
        RECT 0.570 1.130 0.740 1.950 ;
        RECT 1.250 1.300 1.610 1.630 ;
        RECT 0.115 0.960 0.740 1.130 ;
        RECT 1.440 1.030 1.610 1.300 ;
        RECT 1.780 1.290 2.045 2.320 ;
        RECT 2.295 2.200 2.625 2.980 ;
        RECT 2.795 2.370 3.125 3.245 ;
        RECT 3.295 2.200 3.625 2.980 ;
        RECT 3.815 2.290 4.145 3.245 ;
        RECT 2.215 2.030 3.625 2.200 ;
        RECT 4.315 2.120 4.645 2.980 ;
        RECT 2.215 1.030 2.385 2.030 ;
        RECT 4.060 1.950 4.645 2.120 ;
        RECT 0.115 0.350 0.365 0.960 ;
        RECT 1.440 0.860 2.385 1.030 ;
        RECT 0.545 0.085 0.875 0.790 ;
        RECT 1.820 0.350 2.385 0.860 ;
        RECT 2.555 1.020 2.845 1.790 ;
        RECT 4.060 1.030 4.230 1.950 ;
        RECT 4.060 1.020 4.685 1.030 ;
        RECT 2.555 0.850 4.685 1.020 ;
        RECT 3.720 0.085 4.110 0.680 ;
        RECT 4.355 0.440 4.685 0.850 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__and4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hs__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.550 1.780 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 4.825 1.180 5.155 1.590 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.310 1.420 2.755 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.420 3.255 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.050 5.275 1.280 ;
        RECT 0.005 0.245 5.275 1.050 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.835 1.840 4.195 2.980 ;
        RECT 4.025 1.170 4.195 1.840 ;
        RECT 3.815 0.920 4.195 1.170 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.210 2.120 0.540 2.820 ;
        RECT 0.780 2.290 1.110 3.245 ;
        RECT 1.430 2.120 1.760 2.980 ;
        RECT 2.065 2.290 2.395 3.245 ;
        RECT 2.610 2.120 2.940 2.980 ;
        RECT 3.200 2.290 3.530 3.245 ;
        RECT 0.210 1.950 0.935 2.120 ;
        RECT 0.765 1.670 0.935 1.950 ;
        RECT 1.430 1.950 3.665 2.120 ;
        RECT 4.365 2.100 4.615 3.245 ;
        RECT 1.430 1.940 1.760 1.950 ;
        RECT 0.765 1.340 1.260 1.670 ;
        RECT 0.765 1.280 0.935 1.340 ;
        RECT 0.115 1.110 0.935 1.280 ;
        RECT 1.430 1.170 1.600 1.940 ;
        RECT 3.495 1.670 3.665 1.950 ;
        RECT 4.820 1.930 5.165 2.700 ;
        RECT 4.365 1.760 5.165 1.930 ;
        RECT 0.115 0.350 0.365 1.110 ;
        RECT 0.545 0.085 0.875 0.940 ;
        RECT 1.105 0.390 1.600 1.170 ;
        RECT 1.770 1.170 2.100 1.590 ;
        RECT 3.495 1.340 3.855 1.670 ;
        RECT 1.770 1.000 3.645 1.170 ;
        RECT 2.975 0.085 3.305 0.830 ;
        RECT 3.475 0.750 3.645 1.000 ;
        RECT 4.365 0.750 4.535 1.760 ;
        RECT 4.835 0.750 5.165 1.010 ;
        RECT 3.475 0.580 5.165 0.750 ;
        RECT 4.325 0.085 4.655 0.410 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__and4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hs__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.450 1.335 1.780 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.835 1.780 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.965 1.450 6.115 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.350 6.875 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.930 1.455 4.270 1.470 ;
        RECT 1.930 1.240 5.760 1.455 ;
        RECT 1.930 1.140 9.115 1.240 ;
        RECT 0.005 0.245 9.115 1.140 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.760 9.310 3.520 ;
        RECT -0.190 1.660 1.720 1.760 ;
        RECT 5.970 1.660 9.310 1.760 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 7.405 2.150 7.575 2.980 ;
        RECT 7.405 1.820 8.995 2.150 ;
        RECT 8.765 1.150 8.995 1.820 ;
        RECT 7.240 0.980 8.995 1.150 ;
        RECT 7.240 0.350 7.570 0.980 ;
        RECT 8.240 0.770 8.995 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.615 2.290 0.945 3.245 ;
        RECT 1.115 2.460 1.445 2.980 ;
        RECT 1.890 2.630 2.225 3.245 ;
        RECT 1.115 2.290 2.260 2.460 ;
        RECT 0.115 1.950 1.675 2.120 ;
        RECT 1.505 1.280 1.675 1.950 ;
        RECT 1.930 1.450 2.260 2.290 ;
        RECT 2.430 1.765 2.760 2.960 ;
        RECT 2.965 1.935 3.295 3.245 ;
        RECT 3.465 1.765 3.795 2.960 ;
        RECT 3.965 1.935 4.295 3.245 ;
        RECT 4.465 2.120 4.795 2.960 ;
        RECT 4.965 2.290 6.165 3.245 ;
        RECT 6.335 2.120 6.665 2.860 ;
        RECT 6.875 2.290 7.205 3.245 ;
        RECT 7.775 2.320 8.105 3.245 ;
        RECT 8.675 2.320 9.005 3.245 ;
        RECT 4.465 1.950 7.235 2.120 ;
        RECT 4.465 1.765 4.795 1.950 ;
        RECT 2.430 1.595 4.795 1.765 ;
        RECT 7.065 1.650 7.235 1.950 ;
        RECT 2.540 1.360 2.760 1.595 ;
        RECT 0.115 1.110 1.870 1.280 ;
        RECT 0.115 0.350 0.365 1.110 ;
        RECT 0.545 0.085 0.875 0.940 ;
        RECT 1.045 0.585 1.530 0.940 ;
        RECT 1.700 0.925 1.870 1.110 ;
        RECT 2.040 1.095 2.370 1.280 ;
        RECT 2.540 1.095 2.870 1.360 ;
        RECT 3.050 1.255 4.160 1.425 ;
        RECT 2.200 0.925 2.370 1.095 ;
        RECT 3.050 0.925 3.220 1.255 ;
        RECT 3.830 1.095 4.160 1.255 ;
        RECT 4.390 1.280 4.720 1.345 ;
        RECT 7.065 1.320 8.565 1.650 ;
        RECT 4.390 1.180 5.650 1.280 ;
        RECT 4.390 1.110 6.560 1.180 ;
        RECT 4.390 1.095 4.720 1.110 ;
        RECT 1.700 0.755 2.030 0.925 ;
        RECT 2.200 0.755 3.220 0.925 ;
        RECT 3.400 0.925 3.650 1.085 ;
        RECT 5.400 1.010 6.560 1.110 ;
        RECT 4.890 0.925 5.220 0.940 ;
        RECT 3.400 0.755 5.220 0.925 ;
        RECT 1.860 0.585 2.030 0.755 ;
        RECT 4.890 0.665 5.220 0.755 ;
        RECT 5.400 0.665 5.650 1.010 ;
        RECT 1.045 0.255 1.690 0.585 ;
        RECT 1.860 0.255 3.605 0.585 ;
        RECT 5.880 0.085 6.130 0.840 ;
        RECT 6.310 0.450 6.560 1.010 ;
        RECT 6.740 0.085 7.070 1.130 ;
        RECT 7.740 0.085 8.070 0.810 ;
        RECT 8.670 0.085 9.005 0.600 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__and4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hs__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.910 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 1.915 1.240 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 1.470 1.820 1.830 2.980 ;
        RECT 1.660 1.130 1.830 1.820 ;
        RECT 1.475 0.350 1.830 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.470 2.120 0.800 2.980 ;
        RECT 0.970 2.290 1.300 3.245 ;
        RECT 0.470 1.950 1.300 2.120 ;
        RECT 1.130 1.630 1.300 1.950 ;
        RECT 1.130 1.300 1.490 1.630 ;
        RECT 1.130 1.280 1.300 1.300 ;
        RECT 0.115 1.110 1.300 1.280 ;
        RECT 0.115 0.800 0.795 1.110 ;
        RECT 0.975 0.085 1.305 0.940 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__buf_1

#--------EOF---------

MACRO sky130_fd_sc_hs__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.825 1.350 2.275 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.405 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.180 1.315 2.150 ;
        RECT 0.945 0.350 1.275 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.115 2.735 0.825 3.245 ;
        RECT 0.115 1.820 0.420 2.735 ;
        RECT 1.395 2.660 1.725 3.245 ;
        RECT 1.930 2.490 2.285 2.880 ;
        RECT 0.605 2.320 2.285 2.490 ;
        RECT 0.605 1.630 0.775 2.320 ;
        RECT 0.105 1.300 0.775 1.630 ;
        RECT 1.485 1.180 1.655 2.320 ;
        RECT 1.930 1.950 2.285 2.320 ;
        RECT 0.515 0.085 0.765 1.130 ;
        RECT 1.485 1.010 2.285 1.180 ;
        RECT 1.445 0.085 1.775 0.840 ;
        RECT 1.955 0.450 2.285 1.010 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__buf_2

#--------EOF---------

MACRO sky130_fd_sc_hs__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 2.905 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.660 1.970 0.835 2.980 ;
        RECT 1.560 1.970 1.730 2.980 ;
        RECT 0.660 1.800 1.730 1.970 ;
        RECT 0.660 1.410 0.835 1.800 ;
        RECT 0.605 1.180 0.835 1.410 ;
        RECT 0.615 1.130 0.835 1.180 ;
        RECT 0.615 0.960 1.945 1.130 ;
        RECT 0.615 0.350 0.945 0.960 ;
        RECT 1.615 0.350 1.945 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.130 1.820 0.460 3.245 ;
        RECT 1.030 2.140 1.360 3.245 ;
        RECT 1.930 1.820 2.260 3.245 ;
        RECT 2.915 2.370 3.245 3.245 ;
        RECT 2.465 1.950 3.245 2.200 ;
        RECT 1.060 1.300 2.285 1.630 ;
        RECT 2.115 1.130 2.285 1.300 ;
        RECT 3.075 1.130 3.245 1.950 ;
        RECT 0.115 0.085 0.445 1.010 ;
        RECT 2.115 0.960 3.245 1.130 ;
        RECT 1.115 0.085 1.445 0.790 ;
        RECT 2.115 0.085 2.745 0.680 ;
        RECT 2.915 0.350 3.245 0.960 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__buf_4

#--------EOF---------

MACRO sky130_fd_sc_hs__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.837000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.430 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.249300 ;
    PORT
      LAYER li1 ;
        RECT 1.970 1.970 2.300 2.980 ;
        RECT 2.920 1.970 3.250 2.980 ;
        RECT 3.870 1.970 4.200 2.980 ;
        RECT 4.820 1.970 5.155 2.980 ;
        RECT 1.970 1.800 5.155 1.970 ;
        RECT 4.975 1.130 5.145 1.800 ;
        RECT 1.960 0.960 5.145 1.130 ;
        RECT 1.960 0.350 2.130 0.960 ;
        RECT 2.810 0.350 3.140 0.960 ;
        RECT 3.810 0.350 4.140 0.960 ;
        RECT 4.810 0.350 5.145 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.120 2.120 0.450 2.980 ;
        RECT 0.650 2.290 0.820 3.245 ;
        RECT 1.020 2.120 1.350 2.980 ;
        RECT 1.550 2.290 1.800 3.245 ;
        RECT 2.500 2.140 2.750 3.245 ;
        RECT 3.450 2.140 3.700 3.245 ;
        RECT 4.400 2.140 4.650 3.245 ;
        RECT 0.120 1.950 1.770 2.120 ;
        RECT 1.600 1.630 1.770 1.950 ;
        RECT 5.350 1.820 5.600 3.245 ;
        RECT 1.600 1.300 4.805 1.630 ;
        RECT 1.600 1.180 1.770 1.300 ;
        RECT 0.115 1.010 1.770 1.180 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.100 0.350 1.270 1.010 ;
        RECT 1.450 0.085 1.780 0.840 ;
        RECT 2.310 0.085 2.640 0.790 ;
        RECT 3.310 0.085 3.640 0.790 ;
        RECT 4.310 0.085 4.640 0.790 ;
        RECT 5.315 0.085 5.645 1.130 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__buf_8

#--------EOF---------

MACRO sky130_fd_sc_hs__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.674000 ;
    PORT
      LAYER li1 ;
        RECT 7.775 1.350 10.435 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.560 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 10.555 1.240 ;
        RECT 0.000 0.000 10.560 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.750 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.560 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.345600 ;
    PORT
      LAYER met1 ;
        RECT 0.575 1.920 7.255 2.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.560 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 0.130 0.085 0.380 1.130 ;
        RECT 0.560 0.350 0.815 2.980 ;
        RECT 1.095 1.965 1.265 3.245 ;
        RECT 0.985 1.300 1.295 1.780 ;
        RECT 0.990 0.085 1.285 1.130 ;
        RECT 1.465 0.350 1.720 2.980 ;
        RECT 1.965 1.965 2.215 3.245 ;
        RECT 1.890 1.300 2.175 1.780 ;
        RECT 2.415 1.355 2.675 2.980 ;
        RECT 2.945 1.965 3.115 3.245 ;
        RECT 3.310 1.820 3.565 2.980 ;
        RECT 3.845 1.965 4.015 3.245 ;
        RECT 4.215 1.900 4.545 2.980 ;
        RECT 4.745 1.965 4.915 3.245 ;
        RECT 2.345 1.185 2.675 1.355 ;
        RECT 2.845 1.300 3.140 1.780 ;
        RECT 1.895 0.085 2.100 1.130 ;
        RECT 2.345 0.350 2.610 1.185 ;
        RECT 3.310 1.130 3.480 1.820 ;
        RECT 3.735 1.655 4.045 1.780 ;
        RECT 3.655 1.300 4.045 1.655 ;
        RECT 4.215 1.130 4.385 1.900 ;
        RECT 4.675 1.730 4.865 1.780 ;
        RECT 4.555 1.300 4.865 1.730 ;
        RECT 5.115 1.375 5.410 2.980 ;
        RECT 5.645 1.965 5.815 3.245 ;
        RECT 5.035 1.205 5.410 1.375 ;
        RECT 5.580 1.300 5.890 1.780 ;
        RECT 2.790 0.085 2.960 1.015 ;
        RECT 3.220 0.350 3.480 1.130 ;
        RECT 3.650 0.085 3.820 1.130 ;
        RECT 4.000 0.350 4.385 1.130 ;
        RECT 4.555 0.085 4.830 1.130 ;
        RECT 5.035 0.350 5.330 1.205 ;
        RECT 6.060 1.130 6.330 2.980 ;
        RECT 6.545 1.965 6.715 3.245 ;
        RECT 6.500 1.300 6.810 1.780 ;
        RECT 6.980 1.250 7.245 2.980 ;
        RECT 7.445 2.290 7.695 3.245 ;
        RECT 7.865 2.120 8.195 2.980 ;
        RECT 8.395 2.290 8.565 3.245 ;
        RECT 8.765 2.120 9.095 2.980 ;
        RECT 9.295 2.290 9.465 3.245 ;
        RECT 9.665 2.120 9.995 2.980 ;
        RECT 7.420 1.950 9.995 2.120 ;
        RECT 10.195 1.950 10.445 3.245 ;
        RECT 5.500 0.085 5.830 1.035 ;
        RECT 6.000 0.350 6.330 1.130 ;
        RECT 6.500 0.085 6.830 1.130 ;
        RECT 7.000 0.350 7.250 1.250 ;
        RECT 7.420 1.180 7.590 1.950 ;
        RECT 7.420 1.010 9.945 1.180 ;
        RECT 7.430 0.085 7.760 0.840 ;
        RECT 7.940 0.350 8.110 1.010 ;
        RECT 8.290 0.085 8.620 0.840 ;
        RECT 8.800 0.350 8.970 1.010 ;
        RECT 9.150 0.085 9.480 0.840 ;
        RECT 9.695 0.350 9.945 1.010 ;
        RECT 10.115 0.085 10.445 1.130 ;
        RECT 0.000 -0.085 10.560 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 0.635 1.950 0.805 2.120 ;
        RECT 1.515 1.950 1.685 2.120 ;
        RECT 1.055 1.580 1.225 1.750 ;
        RECT 2.470 1.950 2.640 2.120 ;
        RECT 1.950 1.580 2.120 1.750 ;
        RECT 3.360 1.950 3.530 2.120 ;
        RECT 4.300 1.950 4.470 2.120 ;
        RECT 5.195 1.950 5.365 2.120 ;
        RECT 2.910 1.580 3.080 1.750 ;
        RECT 3.800 1.580 3.970 1.750 ;
        RECT 4.680 1.580 4.850 1.750 ;
        RECT 6.095 1.950 6.265 2.120 ;
        RECT 5.650 1.580 5.820 1.750 ;
        RECT 7.025 1.950 7.195 2.120 ;
        RECT 6.565 1.580 6.735 1.750 ;
        RECT 7.420 1.580 7.590 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
      LAYER met1 ;
        RECT 0.985 1.550 7.650 1.780 ;
  END
END sky130_fd_sc_hs__buf_16

#--------EOF---------

MACRO sky130_fd_sc_hs__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__bufbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.570 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.210 7.090 1.240 ;
        RECT 0.005 0.245 7.195 1.210 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.273200 ;
    PORT
      LAYER li1 ;
        RECT 3.565 1.970 3.830 2.980 ;
        RECT 4.495 1.970 4.745 2.980 ;
        RECT 5.385 1.970 5.655 2.980 ;
        RECT 6.285 1.970 6.555 2.980 ;
        RECT 3.565 1.800 6.555 1.970 ;
        RECT 6.255 1.780 6.555 1.800 ;
        RECT 6.255 1.270 7.075 1.780 ;
        RECT 6.255 1.130 6.585 1.270 ;
        RECT 3.475 0.880 6.585 1.130 ;
        RECT 3.475 0.350 3.805 0.880 ;
        RECT 6.255 0.350 6.585 0.880 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.115 2.200 0.380 2.700 ;
        RECT 0.565 2.370 0.920 3.245 ;
        RECT 0.115 1.950 0.920 2.200 ;
        RECT 0.750 1.630 0.920 1.950 ;
        RECT 1.090 1.820 1.480 2.980 ;
        RECT 1.650 1.990 1.980 2.980 ;
        RECT 2.150 2.160 2.380 3.245 ;
        RECT 2.550 1.990 2.880 2.980 ;
        RECT 1.650 1.820 2.880 1.990 ;
        RECT 3.050 1.820 3.380 3.245 ;
        RECT 4.035 2.140 4.290 3.245 ;
        RECT 4.930 2.140 5.205 3.245 ;
        RECT 5.835 2.140 6.105 3.245 ;
        RECT 6.735 1.950 7.040 3.245 ;
        RECT 1.310 1.630 1.480 1.820 ;
        RECT 2.670 1.630 2.880 1.820 ;
        RECT 0.750 1.300 1.140 1.630 ;
        RECT 1.310 1.300 2.500 1.630 ;
        RECT 2.670 1.300 6.020 1.630 ;
        RECT 0.750 1.180 0.920 1.300 ;
        RECT 0.115 1.010 0.920 1.180 ;
        RECT 1.310 1.130 1.480 1.300 ;
        RECT 2.670 1.130 3.125 1.300 ;
        RECT 0.115 0.540 0.445 1.010 ;
        RECT 0.625 0.085 0.955 0.840 ;
        RECT 1.125 0.350 1.480 1.130 ;
        RECT 1.685 0.880 3.125 1.130 ;
        RECT 1.685 0.350 1.935 0.880 ;
        RECT 2.115 0.085 2.445 0.710 ;
        RECT 2.975 0.085 3.305 0.710 ;
        RECT 3.975 0.085 4.305 0.710 ;
        RECT 4.835 0.085 5.165 0.710 ;
        RECT 5.755 0.085 6.085 0.710 ;
        RECT 6.755 0.085 7.085 1.100 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__bufbuf_8

#--------EOF---------

MACRO sky130_fd_sc_hs__bufbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__bufbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.505 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 12.955 1.240 ;
        RECT 0.000 0.000 12.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.150 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.960 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.401600 ;
    PORT
      LAYER met1 ;
        RECT 5.700 1.920 12.380 2.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.645 2.290 0.815 3.245 ;
        RECT 0.115 1.950 0.845 2.120 ;
        RECT 0.675 1.630 0.845 1.950 ;
        RECT 1.015 1.970 1.345 2.980 ;
        RECT 1.545 2.140 1.715 3.245 ;
        RECT 1.915 1.970 2.245 2.980 ;
        RECT 1.015 1.800 2.245 1.970 ;
        RECT 2.490 1.820 2.740 3.245 ;
        RECT 2.940 1.990 3.270 2.980 ;
        RECT 3.470 2.160 3.640 3.245 ;
        RECT 3.840 1.990 4.170 2.980 ;
        RECT 4.370 2.160 4.540 3.245 ;
        RECT 4.750 1.990 5.080 2.980 ;
        RECT 2.940 1.820 5.080 1.990 ;
        RECT 5.280 1.925 5.450 3.245 ;
        RECT 5.660 1.920 5.990 2.980 ;
        RECT 6.160 1.925 6.410 3.245 ;
        RECT 6.610 1.920 6.940 2.980 ;
        RECT 7.140 1.925 7.310 3.245 ;
        RECT 7.510 1.920 7.840 2.980 ;
        RECT 8.040 1.925 8.210 3.245 ;
        RECT 8.410 1.920 8.740 2.980 ;
        RECT 8.940 1.925 9.110 3.245 ;
        RECT 9.310 1.920 9.640 2.980 ;
        RECT 9.840 1.925 10.010 3.245 ;
        RECT 10.210 1.920 10.540 2.980 ;
        RECT 10.740 1.925 10.910 3.245 ;
        RECT 11.110 1.920 11.440 2.980 ;
        RECT 11.640 1.925 11.890 3.245 ;
        RECT 12.060 2.020 12.390 2.980 ;
        RECT 5.660 1.900 5.885 1.920 ;
        RECT 2.045 1.650 2.245 1.800 ;
        RECT 4.845 1.755 5.080 1.820 ;
        RECT 0.675 1.300 1.875 1.630 ;
        RECT 2.045 1.320 4.480 1.650 ;
        RECT 4.845 1.320 5.405 1.755 ;
        RECT 0.675 1.130 0.845 1.300 ;
        RECT 2.045 1.130 2.215 1.320 ;
        RECT 4.845 1.150 5.105 1.320 ;
        RECT 0.130 0.960 0.845 1.130 ;
        RECT 1.070 0.960 2.215 1.130 ;
        RECT 0.130 0.350 0.380 0.960 ;
        RECT 0.560 0.085 0.890 0.790 ;
        RECT 1.070 0.350 1.240 0.960 ;
        RECT 1.420 0.085 1.670 0.790 ;
        RECT 1.855 0.350 2.215 0.960 ;
        RECT 2.415 0.085 2.745 1.130 ;
        RECT 2.915 0.980 5.105 1.150 ;
        RECT 2.915 0.350 3.165 0.980 ;
        RECT 3.345 0.085 3.675 0.810 ;
        RECT 3.845 0.350 4.095 0.980 ;
        RECT 4.275 0.085 4.605 0.810 ;
        RECT 4.775 0.350 5.025 0.980 ;
        RECT 5.275 0.085 5.455 1.130 ;
        RECT 5.635 0.350 5.885 1.900 ;
        RECT 6.055 1.320 6.365 1.750 ;
        RECT 6.610 1.650 6.780 1.920 ;
        RECT 6.065 0.085 6.315 1.130 ;
        RECT 6.535 0.350 6.780 1.650 ;
        RECT 6.950 1.320 7.215 1.750 ;
        RECT 7.510 1.650 7.680 1.920 ;
        RECT 6.960 0.085 7.175 1.130 ;
        RECT 7.385 0.350 7.680 1.650 ;
        RECT 7.850 1.320 8.115 1.750 ;
        RECT 8.410 1.650 8.580 1.920 ;
        RECT 7.850 0.085 8.115 1.130 ;
        RECT 8.285 0.350 8.580 1.650 ;
        RECT 8.750 1.320 9.045 1.750 ;
        RECT 9.310 1.650 9.480 1.920 ;
        RECT 8.750 0.085 9.045 1.130 ;
        RECT 9.215 0.350 9.480 1.650 ;
        RECT 9.650 1.320 9.975 1.750 ;
        RECT 10.210 1.650 10.395 1.920 ;
        RECT 9.665 0.085 9.975 1.130 ;
        RECT 10.145 0.350 10.395 1.650 ;
        RECT 10.565 1.320 10.940 1.750 ;
        RECT 10.575 0.085 10.905 1.130 ;
        RECT 11.110 0.350 11.325 1.920 ;
        RECT 11.495 1.320 11.890 1.750 ;
        RECT 12.060 1.150 12.345 2.020 ;
        RECT 12.590 1.820 12.840 3.245 ;
        RECT 11.505 0.085 11.835 1.130 ;
        RECT 12.015 0.350 12.345 1.150 ;
        RECT 12.515 0.085 12.845 1.130 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 5.760 1.950 5.930 2.120 ;
        RECT 6.675 1.950 6.845 2.120 ;
        RECT 7.595 1.950 7.765 2.120 ;
        RECT 8.485 1.950 8.655 2.120 ;
        RECT 9.405 1.950 9.575 2.120 ;
        RECT 10.295 1.950 10.465 2.120 ;
        RECT 11.195 1.950 11.365 2.120 ;
        RECT 12.115 1.950 12.285 2.120 ;
        RECT 5.180 1.580 5.350 1.750 ;
        RECT 6.125 1.580 6.295 1.750 ;
        RECT 7.000 1.580 7.170 1.750 ;
        RECT 7.900 1.580 8.070 1.750 ;
        RECT 8.820 1.580 8.990 1.750 ;
        RECT 9.730 1.580 9.900 1.750 ;
        RECT 10.675 1.580 10.845 1.750 ;
        RECT 11.600 1.580 11.770 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
      LAYER met1 ;
        RECT 5.110 1.550 11.830 1.780 ;
  END
END sky130_fd_sc_hs__bufbuf_16

#--------EOF---------

MACRO sky130_fd_sc_hs__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__bufinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 6.235 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.385000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.800 4.225 2.070 ;
        RECT 1.060 1.130 1.390 1.800 ;
        RECT 1.060 0.960 4.250 1.130 ;
        RECT 1.060 0.880 3.250 0.960 ;
        RECT 1.060 0.350 1.390 0.880 ;
        RECT 2.060 0.350 2.250 0.880 ;
        RECT 2.920 0.350 3.250 0.880 ;
        RECT 3.920 0.350 4.250 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.115 2.410 0.445 2.980 ;
        RECT 0.615 2.580 0.945 3.245 ;
        RECT 1.515 2.580 1.845 3.245 ;
        RECT 2.415 2.580 2.745 3.245 ;
        RECT 3.315 2.580 3.645 3.245 ;
        RECT 4.345 2.580 4.675 3.245 ;
        RECT 0.115 2.240 4.565 2.410 ;
        RECT 0.115 1.950 0.445 2.240 ;
        RECT 0.720 1.180 0.890 2.240 ;
        RECT 4.395 1.970 4.565 2.240 ;
        RECT 4.845 2.310 5.175 2.980 ;
        RECT 5.345 2.480 5.675 3.245 ;
        RECT 5.845 2.310 6.125 2.980 ;
        RECT 4.845 2.140 6.125 2.310 ;
        RECT 4.395 1.800 5.605 1.970 ;
        RECT 1.665 1.300 4.820 1.630 ;
        RECT 4.990 1.320 5.605 1.800 ;
        RECT 0.130 1.010 0.890 1.180 ;
        RECT 4.650 1.130 4.820 1.300 ;
        RECT 5.795 1.130 6.125 2.140 ;
        RECT 0.130 0.350 0.380 1.010 ;
        RECT 4.650 0.880 6.125 1.130 ;
        RECT 0.560 0.085 0.890 0.840 ;
        RECT 1.560 0.085 1.890 0.710 ;
        RECT 2.420 0.085 2.750 0.710 ;
        RECT 3.420 0.085 3.750 0.790 ;
        RECT 4.420 0.085 4.750 0.710 ;
        RECT 4.920 0.350 5.125 0.880 ;
        RECT 5.295 0.085 5.625 0.710 ;
        RECT 5.795 0.350 6.125 0.880 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__bufinv_8

#--------EOF---------

MACRO sky130_fd_sc_hs__bufinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__bufinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.837000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.430 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.000 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 11.995 1.240 ;
        RECT 0.000 0.000 12.000 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 12.190 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.000 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.390400 ;
    PORT
      LAYER met1 ;
        RECT 4.660 1.920 11.400 2.150 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.000 3.415 ;
        RECT 0.120 2.120 0.450 2.980 ;
        RECT 0.650 2.290 0.820 3.245 ;
        RECT 1.020 2.120 1.350 2.980 ;
        RECT 1.550 2.290 1.720 3.245 ;
        RECT 0.120 1.950 1.770 2.120 ;
        RECT 1.600 1.630 1.770 1.950 ;
        RECT 1.940 1.970 2.270 2.980 ;
        RECT 2.470 2.140 2.640 3.245 ;
        RECT 2.840 1.970 3.170 2.980 ;
        RECT 3.370 2.140 3.540 3.245 ;
        RECT 3.740 1.970 4.070 2.980 ;
        RECT 1.940 1.800 4.070 1.970 ;
        RECT 4.270 1.920 4.440 3.245 ;
        RECT 4.640 2.020 4.970 2.980 ;
        RECT 4.615 1.920 4.970 2.020 ;
        RECT 5.170 1.920 5.340 3.245 ;
        RECT 5.540 2.020 5.870 2.980 ;
        RECT 5.510 1.920 5.870 2.020 ;
        RECT 6.070 1.920 6.240 3.245 ;
        RECT 6.440 2.020 6.770 2.980 ;
        RECT 6.420 1.920 6.770 2.020 ;
        RECT 6.970 1.920 7.140 3.245 ;
        RECT 7.340 1.920 7.670 2.980 ;
        RECT 7.870 1.920 8.040 3.245 ;
        RECT 8.240 2.020 8.570 2.980 ;
        RECT 8.265 1.920 8.570 2.020 ;
        RECT 8.770 1.920 8.995 3.245 ;
        RECT 9.190 2.020 9.520 2.980 ;
        RECT 9.195 1.920 9.520 2.020 ;
        RECT 9.720 1.920 9.955 3.245 ;
        RECT 10.140 2.020 10.470 2.980 ;
        RECT 10.125 1.920 10.470 2.020 ;
        RECT 10.670 1.920 10.885 3.245 ;
        RECT 11.090 2.020 11.420 2.980 ;
        RECT 3.740 1.750 4.070 1.800 ;
        RECT 1.600 1.300 3.460 1.630 ;
        RECT 3.740 1.300 4.435 1.750 ;
        RECT 1.600 1.180 1.770 1.300 ;
        RECT 0.115 1.010 1.770 1.180 ;
        RECT 3.685 1.130 3.935 1.300 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.115 0.350 1.285 1.010 ;
        RECT 1.975 0.960 3.935 1.130 ;
        RECT 1.465 0.085 1.795 0.840 ;
        RECT 1.975 0.350 2.145 0.960 ;
        RECT 2.325 0.085 2.575 0.790 ;
        RECT 2.755 0.350 3.005 0.960 ;
        RECT 3.185 0.085 3.515 0.790 ;
        RECT 3.685 0.350 3.935 0.960 ;
        RECT 4.115 0.085 4.445 1.130 ;
        RECT 4.615 0.350 4.865 1.920 ;
        RECT 5.035 1.300 5.305 1.750 ;
        RECT 5.045 0.085 5.295 1.105 ;
        RECT 5.510 0.350 5.725 1.920 ;
        RECT 5.900 1.300 6.230 1.750 ;
        RECT 5.905 0.085 6.235 1.105 ;
        RECT 6.420 0.350 6.655 1.920 ;
        RECT 6.840 1.300 7.170 1.750 ;
        RECT 6.835 0.085 7.165 1.105 ;
        RECT 7.340 0.350 7.585 1.920 ;
        RECT 7.760 1.300 8.090 1.750 ;
        RECT 7.765 0.085 8.095 1.105 ;
        RECT 8.265 0.350 8.515 1.920 ;
        RECT 8.685 1.300 9.015 1.750 ;
        RECT 8.695 0.085 9.025 1.105 ;
        RECT 9.195 0.350 9.445 1.920 ;
        RECT 9.615 1.300 9.945 1.750 ;
        RECT 9.625 0.085 9.955 1.105 ;
        RECT 10.125 0.350 10.375 1.920 ;
        RECT 11.055 1.790 11.420 2.020 ;
        RECT 11.620 1.820 11.870 3.245 ;
        RECT 10.545 1.300 10.875 1.750 ;
        RECT 10.555 0.085 10.885 1.105 ;
        RECT 11.055 0.350 11.385 1.790 ;
        RECT 11.555 0.085 11.885 1.130 ;
        RECT 0.000 -0.085 12.000 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 4.730 1.950 4.900 2.120 ;
        RECT 5.620 1.950 5.790 2.120 ;
        RECT 6.520 1.950 6.690 2.120 ;
        RECT 7.420 1.950 7.590 2.120 ;
        RECT 8.320 1.950 8.490 2.120 ;
        RECT 9.270 1.950 9.440 2.120 ;
        RECT 10.220 1.950 10.390 2.120 ;
        RECT 11.170 1.950 11.340 2.120 ;
        RECT 4.225 1.580 4.395 1.750 ;
        RECT 5.090 1.580 5.260 1.750 ;
        RECT 5.980 1.580 6.150 1.750 ;
        RECT 6.920 1.580 7.090 1.750 ;
        RECT 7.835 1.580 8.005 1.750 ;
        RECT 8.765 1.580 8.935 1.750 ;
        RECT 9.690 1.580 9.860 1.750 ;
        RECT 10.625 1.580 10.795 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
      LAYER met1 ;
        RECT 4.155 1.550 10.855 1.780 ;
  END
END sky130_fd_sc_hs__bufinv_16

#--------EOF---------

MACRO sky130_fd_sc_hs__clkbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.835 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.900 1.880 0.920 ;
        RECT 0.005 0.245 1.915 0.900 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449400 ;
    PORT
      LAYER li1 ;
        RECT 1.345 1.820 1.805 2.980 ;
        RECT 1.565 0.790 1.805 1.820 ;
        RECT 1.475 0.350 1.805 0.790 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.345 2.120 0.675 2.980 ;
        RECT 0.845 2.290 1.175 3.245 ;
        RECT 0.345 1.950 1.175 2.120 ;
        RECT 1.005 1.630 1.175 1.950 ;
        RECT 1.005 1.130 1.395 1.630 ;
        RECT 0.115 0.960 1.395 1.130 ;
        RECT 0.115 0.350 0.445 0.960 ;
        RECT 0.615 0.085 1.305 0.680 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__clkbuf_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.010 1.495 2.150 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 1.915 0.920 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453600 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.820 0.885 2.150 ;
        RECT 0.715 0.790 0.885 1.820 ;
        RECT 0.545 0.350 0.885 0.790 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.105 2.660 0.435 3.245 ;
        RECT 1.005 2.660 1.335 3.245 ;
        RECT 1.535 2.490 1.835 2.980 ;
        RECT 0.215 2.320 1.835 2.490 ;
        RECT 0.215 1.630 0.385 2.320 ;
        RECT 0.215 0.960 0.545 1.630 ;
        RECT 1.665 0.810 1.835 2.320 ;
        RECT 0.115 0.085 0.365 0.790 ;
        RECT 1.055 0.085 1.305 0.810 ;
        RECT 1.475 0.350 1.835 0.810 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__clkbuf_2

#--------EOF---------

MACRO sky130_fd_sc_hs__clkbuf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.080 2.455 1.410 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 2.875 0.920 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 2.090 0.815 2.980 ;
        RECT 1.465 2.090 1.795 2.980 ;
        RECT 0.535 1.920 1.795 2.090 ;
        RECT 0.535 1.150 0.705 1.920 ;
        RECT 0.535 0.980 1.750 1.150 ;
        RECT 0.560 0.350 0.890 0.980 ;
        RECT 1.420 0.350 1.750 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.015 2.260 1.265 3.245 ;
        RECT 1.995 1.920 2.245 3.245 ;
        RECT 2.415 1.750 2.795 2.980 ;
        RECT 0.875 1.580 2.795 1.750 ;
        RECT 0.875 1.350 1.885 1.580 ;
        RECT 2.625 0.810 2.795 1.580 ;
        RECT 0.130 0.085 0.380 0.810 ;
        RECT 1.070 0.085 1.240 0.810 ;
        RECT 1.920 0.085 2.250 0.810 ;
        RECT 2.420 0.480 2.795 0.810 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__clkbuf_4

#--------EOF---------

MACRO sky130_fd_sc_hs__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.095 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.275 0.920 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.841700 ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.860 1.880 2.980 ;
        RECT 2.585 1.860 2.845 2.980 ;
        RECT 3.415 1.860 3.680 2.980 ;
        RECT 4.385 1.860 4.645 2.980 ;
        RECT 1.615 1.690 5.155 1.860 ;
        RECT 4.710 1.180 5.155 1.690 ;
        RECT 4.710 1.020 4.880 1.180 ;
        RECT 1.615 0.850 4.880 1.020 ;
        RECT 1.615 0.350 1.945 0.850 ;
        RECT 2.615 0.350 2.865 0.850 ;
        RECT 3.555 0.350 3.725 0.850 ;
        RECT 4.485 0.350 4.655 0.850 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.115 1.950 0.445 3.245 ;
        RECT 0.615 2.120 0.945 2.980 ;
        RECT 1.115 2.290 1.445 3.245 ;
        RECT 0.615 1.950 1.445 2.120 ;
        RECT 2.065 2.030 2.395 3.245 ;
        RECT 3.045 2.030 3.215 3.245 ;
        RECT 3.865 2.030 4.195 3.245 ;
        RECT 4.830 2.030 5.160 3.245 ;
        RECT 1.275 1.520 1.445 1.950 ;
        RECT 1.275 1.190 4.515 1.520 ;
        RECT 1.275 1.150 1.445 1.190 ;
        RECT 0.615 0.980 1.445 1.150 ;
        RECT 0.115 0.085 0.445 0.810 ;
        RECT 0.615 0.350 0.945 0.980 ;
        RECT 1.115 0.085 1.445 0.810 ;
        RECT 2.115 0.085 2.445 0.680 ;
        RECT 3.045 0.085 3.375 0.680 ;
        RECT 3.905 0.085 4.305 0.680 ;
        RECT 4.835 0.085 5.165 0.680 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__clkbuf_8

#--------EOF---------

MACRO sky130_fd_sc_hs__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.795 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 9.595 0.920 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.628800 ;
    PORT
      LAYER met1 ;
        RECT 2.390 1.920 9.090 2.150 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.120 1.950 0.370 3.245 ;
        RECT 0.570 2.120 0.900 2.980 ;
        RECT 1.100 2.290 1.270 3.245 ;
        RECT 1.470 2.120 1.800 2.980 ;
        RECT 2.000 2.290 2.250 3.245 ;
        RECT 2.430 2.120 2.660 2.980 ;
        RECT 0.570 1.950 2.135 2.120 ;
        RECT 1.965 1.410 2.135 1.950 ;
        RECT 1.965 1.180 2.210 1.410 ;
        RECT 1.965 1.150 2.135 1.180 ;
        RECT 0.545 0.980 2.135 1.150 ;
        RECT 0.115 0.085 0.365 0.810 ;
        RECT 0.545 0.350 0.795 0.980 ;
        RECT 0.975 0.085 1.225 0.810 ;
        RECT 1.425 0.350 1.675 0.980 ;
        RECT 1.855 0.085 2.185 0.810 ;
        RECT 2.390 0.350 2.660 2.120 ;
        RECT 2.830 2.030 3.160 3.245 ;
        RECT 3.340 1.860 3.545 2.980 ;
        RECT 3.730 2.030 4.060 3.245 ;
        RECT 4.230 1.860 4.430 2.980 ;
        RECT 4.630 2.030 4.960 3.245 ;
        RECT 5.140 1.860 5.350 2.980 ;
        RECT 5.530 2.030 5.860 3.245 ;
        RECT 6.040 1.860 6.245 2.980 ;
        RECT 6.430 2.030 6.760 3.245 ;
        RECT 6.945 1.860 7.150 2.980 ;
        RECT 7.330 2.030 7.660 3.245 ;
        RECT 7.840 1.860 8.050 2.980 ;
        RECT 8.230 2.030 8.560 3.245 ;
        RECT 8.750 1.860 8.970 2.980 ;
        RECT 9.150 2.030 9.480 3.245 ;
        RECT 3.275 1.690 3.545 1.860 ;
        RECT 4.170 1.690 4.430 1.860 ;
        RECT 5.025 1.690 5.350 1.860 ;
        RECT 5.935 1.690 6.245 1.860 ;
        RECT 6.865 1.690 7.150 1.860 ;
        RECT 7.795 1.690 8.050 1.860 ;
        RECT 8.725 1.830 8.970 1.860 ;
        RECT 2.835 1.190 3.105 1.520 ;
        RECT 2.865 0.085 3.035 0.680 ;
        RECT 3.275 0.350 3.500 1.690 ;
        RECT 3.670 1.190 4.000 1.520 ;
        RECT 4.170 0.745 4.340 1.690 ;
        RECT 4.510 1.190 4.840 1.520 ;
        RECT 3.670 0.085 3.895 0.725 ;
        RECT 4.075 0.350 4.340 0.745 ;
        RECT 4.510 0.085 4.835 0.740 ;
        RECT 5.025 0.350 5.255 1.690 ;
        RECT 5.425 1.190 5.755 1.520 ;
        RECT 5.435 0.085 5.765 0.680 ;
        RECT 5.935 0.350 6.185 1.690 ;
        RECT 6.365 1.190 6.695 1.520 ;
        RECT 6.365 0.085 6.695 0.680 ;
        RECT 6.865 0.350 7.115 1.690 ;
        RECT 7.295 1.190 7.625 1.520 ;
        RECT 7.295 0.085 7.625 0.680 ;
        RECT 7.795 0.350 8.045 1.690 ;
        RECT 8.225 1.190 8.555 1.520 ;
        RECT 8.225 0.085 8.555 0.680 ;
        RECT 8.725 0.350 8.975 1.830 ;
        RECT 9.155 0.085 9.485 0.745 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 2.460 1.950 2.630 2.120 ;
        RECT 2.010 1.210 2.180 1.380 ;
        RECT 3.360 1.950 3.530 2.120 ;
        RECT 4.245 1.950 4.415 2.120 ;
        RECT 5.160 1.950 5.330 2.120 ;
        RECT 6.060 1.950 6.230 2.120 ;
        RECT 6.960 1.950 7.130 2.120 ;
        RECT 7.860 1.950 8.030 2.120 ;
        RECT 8.780 1.950 8.950 2.120 ;
        RECT 2.890 1.210 3.060 1.380 ;
        RECT 3.750 1.210 3.920 1.380 ;
        RECT 4.590 1.210 4.760 1.380 ;
        RECT 5.505 1.210 5.675 1.380 ;
        RECT 6.445 1.210 6.615 1.380 ;
        RECT 7.375 1.210 7.545 1.380 ;
        RECT 8.305 1.210 8.475 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
      LAYER met1 ;
        RECT 1.940 1.180 8.640 1.410 ;
  END
END sky130_fd_sc_hs__clkbuf_16

#--------EOF---------

MACRO sky130_fd_sc_hs__clkdlyinv3sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkdlyinv3sd1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 2.785 0.920 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424900 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.815 2.795 3.060 ;
        RECT 2.530 0.755 2.795 1.815 ;
        RECT 2.435 0.355 2.795 0.755 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.650 1.745 2.900 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.625 1.745 2.650 ;
        RECT 1.935 1.900 2.265 3.245 ;
        RECT 1.475 1.295 2.360 1.625 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.305 1.720 1.295 ;
        RECT 1.935 0.085 2.265 0.750 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__clkdlyinv3sd1_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkdlyinv3sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkdlyinv3sd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 2.785 0.920 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424900 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.815 2.795 3.060 ;
        RECT 2.530 0.755 2.795 1.815 ;
        RECT 2.435 0.355 2.795 0.755 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.650 1.745 2.900 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.625 1.745 2.650 ;
        RECT 1.935 1.900 2.265 3.245 ;
        RECT 1.475 1.295 2.360 1.625 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.305 1.720 1.295 ;
        RECT 1.935 0.085 2.265 0.750 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__clkdlyinv3sd2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkdlyinv3sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkdlyinv3sd3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 2.785 0.920 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424900 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.815 2.795 3.060 ;
        RECT 2.530 0.755 2.795 1.815 ;
        RECT 2.435 0.355 2.795 0.755 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.650 1.745 2.900 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.625 1.745 2.650 ;
        RECT 1.935 1.900 2.265 3.245 ;
        RECT 1.475 1.295 2.360 1.625 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.305 1.720 1.295 ;
        RECT 1.935 0.085 2.265 0.750 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__clkdlyinv3sd3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkdlyinv5sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkdlyinv5sd1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 5.180 0.920 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424900 ;
    PORT
      LAYER li1 ;
        RECT 4.830 1.900 5.190 3.060 ;
        RECT 4.925 0.755 5.190 1.900 ;
        RECT 4.830 0.355 5.190 0.755 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.650 1.745 2.900 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.470 1.745 2.650 ;
        RECT 1.915 1.940 2.265 3.245 ;
        RECT 1.475 1.140 2.510 1.470 ;
        RECT 2.800 1.390 2.970 2.980 ;
        RECT 3.415 1.730 3.655 2.980 ;
        RECT 4.330 1.900 4.660 3.245 ;
        RECT 3.415 1.560 4.755 1.730 ;
        RECT 2.800 1.220 4.005 1.390 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.305 1.720 1.140 ;
        RECT 1.915 0.085 2.265 0.745 ;
        RECT 2.800 0.415 2.970 1.220 ;
        RECT 4.530 1.050 4.755 1.560 ;
        RECT 3.370 0.925 4.755 1.050 ;
        RECT 3.370 0.880 4.700 0.925 ;
        RECT 3.370 0.400 3.700 0.880 ;
        RECT 4.330 0.085 4.660 0.670 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__clkdlyinv5sd1_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkdlyinv5sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkdlyinv5sd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 5.180 0.920 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424900 ;
    PORT
      LAYER li1 ;
        RECT 4.830 1.900 5.190 3.060 ;
        RECT 4.925 0.755 5.190 1.900 ;
        RECT 4.830 0.355 5.190 0.755 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.650 1.745 2.900 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.470 1.745 2.650 ;
        RECT 1.915 1.940 2.265 3.245 ;
        RECT 1.475 1.140 2.510 1.470 ;
        RECT 2.800 1.390 2.970 2.980 ;
        RECT 3.415 1.730 3.655 2.980 ;
        RECT 4.330 1.900 4.660 3.245 ;
        RECT 3.415 1.560 4.755 1.730 ;
        RECT 2.800 1.220 4.005 1.390 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.305 1.720 1.140 ;
        RECT 1.915 0.085 2.265 0.745 ;
        RECT 2.800 0.415 2.970 1.220 ;
        RECT 4.530 1.050 4.755 1.560 ;
        RECT 3.370 0.925 4.755 1.050 ;
        RECT 3.370 0.880 4.700 0.925 ;
        RECT 3.370 0.400 3.700 0.880 ;
        RECT 4.330 0.085 4.660 0.670 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__clkdlyinv5sd2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkdlyinv5sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkdlyinv5sd3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.231000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 5.180 0.920 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424900 ;
    PORT
      LAYER li1 ;
        RECT 4.830 1.900 5.190 3.060 ;
        RECT 4.925 0.755 5.190 1.900 ;
        RECT 4.830 0.355 5.190 0.755 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.650 1.745 2.900 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.470 1.745 2.650 ;
        RECT 1.915 1.940 2.265 3.245 ;
        RECT 1.475 1.140 2.510 1.470 ;
        RECT 2.800 1.390 2.970 2.980 ;
        RECT 3.415 1.730 3.655 2.980 ;
        RECT 4.330 1.900 4.660 3.245 ;
        RECT 3.415 1.560 4.755 1.730 ;
        RECT 2.800 1.220 4.005 1.390 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.305 1.720 1.140 ;
        RECT 1.915 0.085 2.265 0.745 ;
        RECT 2.800 0.415 2.970 1.220 ;
        RECT 4.530 1.050 4.755 1.560 ;
        RECT 3.370 0.925 4.755 1.050 ;
        RECT 3.370 0.880 4.700 0.925 ;
        RECT 3.370 0.400 3.700 0.880 ;
        RECT 4.330 0.085 4.660 0.670 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__clkdlyinv5sd3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkinv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkinv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.315000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.780 0.755 1.930 ;
        RECT 0.125 1.180 0.755 1.780 ;
        RECT 0.425 0.920 0.755 1.180 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.790 1.020 0.920 ;
        RECT 0.005 0.245 1.435 0.790 ;
        RECT 0.000 0.000 1.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.440 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.477350 ;
    PORT
      LAYER li1 ;
        RECT 0.555 2.430 0.835 2.955 ;
        RECT 0.555 2.100 1.325 2.430 ;
        RECT 1.085 0.680 1.325 2.100 ;
        RECT 0.615 0.350 1.325 0.680 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.440 3.415 ;
        RECT 0.105 2.100 0.355 3.245 ;
        RECT 1.005 2.600 1.335 3.245 ;
        RECT 0.115 0.085 0.445 0.750 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
  END
END sky130_fd_sc_hs__clkinv_1

#--------EOF---------

MACRO sky130_fd_sc_hs__clkinv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkinv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.315 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 1.915 0.950 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.994000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 2.120 0.450 2.980 ;
        RECT 1.020 2.120 1.350 2.980 ;
        RECT 0.120 1.950 1.795 2.120 ;
        RECT 1.565 1.180 1.795 1.950 ;
        RECT 0.615 1.010 1.795 1.180 ;
        RECT 0.615 0.510 1.305 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.650 2.290 0.820 3.245 ;
        RECT 1.550 2.290 1.800 3.245 ;
        RECT 0.115 0.085 0.445 0.840 ;
        RECT 1.475 0.085 1.805 0.840 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__clkinv_2

#--------EOF---------

MACRO sky130_fd_sc_hs__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkinv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 2.755 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.355 0.950 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.432200 ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.120 0.895 2.980 ;
        RECT 1.465 2.120 1.795 2.980 ;
        RECT 2.415 2.120 2.745 2.980 ;
        RECT 0.265 1.950 3.235 2.120 ;
        RECT 0.265 1.180 0.435 1.950 ;
        RECT 3.005 1.180 3.235 1.950 ;
        RECT 0.265 1.010 3.235 1.180 ;
        RECT 0.990 0.455 1.745 1.010 ;
        RECT 2.415 0.380 2.745 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.290 0.365 3.245 ;
        RECT 1.095 2.290 1.265 3.245 ;
        RECT 1.995 2.290 2.245 3.245 ;
        RECT 2.915 2.290 3.245 3.245 ;
        RECT 0.115 0.085 0.820 0.710 ;
        RECT 1.915 0.085 2.245 0.840 ;
        RECT 2.915 0.085 3.245 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__clkinv_4

#--------EOF---------

MACRO sky130_fd_sc_hs__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.520000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.350 5.715 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 6.235 0.950 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.242400 ;
    PORT
      LAYER li1 ;
        RECT 0.590 2.120 0.920 2.980 ;
        RECT 1.540 2.120 1.870 2.980 ;
        RECT 2.490 2.120 2.820 2.980 ;
        RECT 3.440 2.120 3.770 2.980 ;
        RECT 4.390 2.120 4.720 2.980 ;
        RECT 5.340 2.120 5.670 2.980 ;
        RECT 0.285 1.950 6.115 2.120 ;
        RECT 0.285 1.180 0.455 1.950 ;
        RECT 5.885 1.180 6.115 1.950 ;
        RECT 0.285 1.010 6.115 1.180 ;
        RECT 0.615 0.460 2.625 1.010 ;
        RECT 3.295 0.445 3.625 1.010 ;
        RECT 4.295 0.445 4.625 1.010 ;
        RECT 5.295 0.445 5.625 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.115 2.290 0.390 3.245 ;
        RECT 1.120 2.290 1.370 3.245 ;
        RECT 2.070 2.290 2.320 3.245 ;
        RECT 3.020 2.290 3.270 3.245 ;
        RECT 3.970 2.290 4.220 3.245 ;
        RECT 4.920 2.290 5.170 3.245 ;
        RECT 5.870 2.290 6.120 3.245 ;
        RECT 0.115 0.085 0.445 0.775 ;
        RECT 2.795 0.085 3.125 0.775 ;
        RECT 3.795 0.085 4.125 0.775 ;
        RECT 4.795 0.085 5.125 0.775 ;
        RECT 5.795 0.085 6.125 0.775 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__clkinv_8

#--------EOF---------

MACRO sky130_fd_sc_hs__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.040000 ;
    PORT
      LAYER met1 ;
        RECT 0.985 1.180 10.935 1.410 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.520 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.820 7.820 0.950 ;
        RECT 0.005 0.245 9.935 0.820 ;
        RECT 0.000 0.000 11.520 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.710 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.520 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.040000 ;
    PORT
      LAYER met1 ;
        RECT 0.575 1.920 10.935 2.150 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.115 1.900 0.445 3.245 ;
        RECT 0.625 1.820 0.815 2.980 ;
        RECT 1.015 1.820 1.265 3.245 ;
        RECT 1.465 1.885 1.795 2.980 ;
        RECT 0.115 0.085 0.445 0.840 ;
        RECT 0.625 0.775 0.805 1.820 ;
        RECT 0.975 1.150 1.295 1.650 ;
        RECT 0.615 0.380 0.805 0.775 ;
        RECT 0.975 0.085 1.260 0.840 ;
        RECT 1.465 0.775 1.695 1.885 ;
        RECT 1.995 1.820 2.165 3.245 ;
        RECT 2.365 1.885 2.695 2.980 ;
        RECT 1.865 1.150 2.195 1.650 ;
        RECT 1.440 0.380 1.700 0.775 ;
        RECT 1.885 0.085 2.165 0.840 ;
        RECT 2.365 0.775 2.665 1.885 ;
        RECT 2.895 1.820 3.065 3.245 ;
        RECT 2.835 1.150 3.165 1.650 ;
        RECT 2.350 0.380 2.665 0.775 ;
        RECT 2.845 0.085 3.095 0.840 ;
        RECT 3.335 0.775 3.595 2.980 ;
        RECT 3.795 1.820 3.965 3.245 ;
        RECT 4.165 1.900 4.495 2.980 ;
        RECT 4.165 1.850 4.525 1.900 ;
        RECT 3.765 1.150 4.095 1.650 ;
        RECT 3.300 0.380 3.595 0.775 ;
        RECT 3.765 0.085 4.095 0.840 ;
        RECT 4.265 0.380 4.525 1.850 ;
        RECT 4.695 1.820 4.865 3.245 ;
        RECT 5.065 2.010 5.395 2.980 ;
        RECT 5.065 1.850 5.425 2.010 ;
        RECT 4.755 1.150 5.085 1.650 ;
        RECT 4.765 0.085 5.085 0.840 ;
        RECT 5.255 0.775 5.425 1.850 ;
        RECT 5.595 1.820 5.845 3.245 ;
        RECT 6.015 1.820 6.330 2.980 ;
        RECT 6.510 1.820 6.795 3.245 ;
        RECT 6.095 1.760 6.330 1.820 ;
        RECT 5.595 1.150 5.925 1.650 ;
        RECT 6.095 1.010 6.340 1.760 ;
        RECT 6.545 1.150 6.875 1.650 ;
        RECT 5.255 0.380 5.525 0.775 ;
        RECT 5.695 0.085 5.980 0.840 ;
        RECT 6.160 0.785 6.340 1.010 ;
        RECT 6.160 0.380 6.385 0.785 ;
        RECT 6.555 0.085 6.875 0.840 ;
        RECT 7.045 0.380 7.290 2.980 ;
        RECT 7.475 1.820 7.805 3.245 ;
        RECT 8.005 1.820 8.175 2.980 ;
        RECT 8.375 1.820 8.625 3.245 ;
        RECT 8.905 1.820 9.075 2.980 ;
        RECT 9.275 1.820 9.605 3.245 ;
        RECT 9.805 1.820 9.975 2.980 ;
        RECT 10.175 1.820 10.505 3.245 ;
        RECT 10.705 1.820 10.875 2.980 ;
        RECT 11.075 1.820 11.405 3.245 ;
        RECT 7.525 1.150 10.915 1.650 ;
        RECT 7.485 0.085 9.825 0.710 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 0.635 1.950 0.805 2.120 ;
        RECT 1.545 1.950 1.715 2.120 ;
        RECT 1.045 1.210 1.215 1.380 ;
        RECT 2.445 1.950 2.615 2.120 ;
        RECT 1.945 1.210 2.115 1.380 ;
        RECT 3.375 1.950 3.545 2.120 ;
        RECT 2.915 1.210 3.085 1.380 ;
        RECT 4.245 1.950 4.415 2.120 ;
        RECT 3.845 1.210 4.015 1.380 ;
        RECT 5.145 1.950 5.315 2.120 ;
        RECT 4.835 1.210 5.005 1.380 ;
        RECT 6.095 1.950 6.265 2.120 ;
        RECT 7.075 1.950 7.245 2.120 ;
        RECT 5.675 1.210 5.845 1.380 ;
        RECT 6.625 1.210 6.795 1.380 ;
        RECT 8.005 1.950 8.175 2.120 ;
        RECT 8.905 1.950 9.075 2.120 ;
        RECT 9.805 1.950 9.975 2.120 ;
        RECT 10.705 1.950 10.875 2.120 ;
        RECT 7.745 1.210 7.915 1.380 ;
        RECT 8.105 1.210 8.275 1.380 ;
        RECT 8.465 1.210 8.635 1.380 ;
        RECT 8.825 1.210 8.995 1.380 ;
        RECT 9.185 1.210 9.355 1.380 ;
        RECT 9.545 1.210 9.715 1.380 ;
        RECT 9.905 1.210 10.075 1.380 ;
        RECT 10.265 1.210 10.435 1.380 ;
        RECT 10.625 1.210 10.795 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
  END
END sky130_fd_sc_hs__clkinv_16

#--------EOF---------

MACRO sky130_fd_sc_hs__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__conb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.000 1.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.440 3.575 ;
    END
  END VPWR
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.845 0.395 2.335 ;
        RECT 0.085 0.255 0.615 0.845 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.825 2.485 1.355 3.075 ;
        RECT 1.055 0.995 1.355 2.485 ;
    END
  END LO
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.440 3.415 ;
        RECT 0.285 2.505 0.615 3.245 ;
        RECT 0.825 0.085 1.155 0.825 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
  END
END sky130_fd_sc_hs__conb_1

#--------EOF---------

MACRO sky130_fd_sc_hs__decap_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.245 1.890 0.975 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.095 1.930 0.425 3.245 ;
        RECT 0.170 0.085 0.740 1.585 ;
        RECT 1.145 1.250 1.715 3.245 ;
        RECT 1.450 0.085 1.780 0.805 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__decap_4

#--------EOF---------

MACRO sky130_fd_sc_hs__decap_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__decap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.245 3.165 0.975 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.095 1.930 0.425 3.245 ;
        RECT 0.170 0.085 0.740 1.585 ;
        RECT 1.145 1.250 2.080 3.245 ;
        RECT 2.660 1.940 2.990 3.245 ;
        RECT 1.450 0.085 1.780 0.805 ;
        RECT 2.355 0.085 3.055 1.580 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__decap_8

#--------EOF---------

MACRO sky130_fd_sc_hs__dfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfbbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.495 1.780 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.925 1.180 2.755 1.510 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.350 11.015 1.780 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER met1 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 8.735 2.105 9.025 2.150 ;
        RECT 5.375 1.965 9.025 2.105 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 8.735 1.920 9.025 1.965 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.205 1.250 6.650 1.275 ;
        RECT 10.465 1.250 11.980 1.295 ;
        RECT 4.205 1.240 11.980 1.250 ;
        RECT 0.005 1.145 1.415 1.240 ;
        RECT 4.205 1.145 13.435 1.240 ;
        RECT 0.005 0.245 13.435 1.145 ;
        RECT 0.000 0.000 13.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.440 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.519000 ;
    PORT
      LAYER li1 ;
        RECT 13.005 0.350 13.340 2.980 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.513400 ;
    PORT
      LAYER li1 ;
        RECT 11.575 1.820 11.925 2.980 ;
        RECT 11.755 1.150 11.925 1.820 ;
        RECT 11.555 0.405 11.925 1.150 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.440 3.415 ;
        RECT 0.105 2.120 0.435 2.980 ;
        RECT 0.635 2.290 0.805 3.245 ;
        RECT 1.005 2.905 2.125 3.075 ;
        RECT 0.105 1.950 0.835 2.120 ;
        RECT 0.665 1.630 0.835 1.950 ;
        RECT 1.005 1.820 1.415 2.905 ;
        RECT 0.665 1.300 1.075 1.630 ;
        RECT 0.665 1.130 0.835 1.300 ;
        RECT 1.245 1.130 1.415 1.820 ;
        RECT 0.115 0.960 0.835 1.130 ;
        RECT 0.115 0.350 0.365 0.960 ;
        RECT 0.545 0.085 0.875 0.790 ;
        RECT 1.055 0.350 1.415 1.130 ;
        RECT 1.585 2.405 1.785 2.735 ;
        RECT 1.585 1.010 1.755 2.405 ;
        RECT 1.955 1.855 2.125 2.905 ;
        RECT 2.295 2.525 2.465 3.245 ;
        RECT 2.635 2.905 4.530 3.075 ;
        RECT 2.635 2.355 2.805 2.905 ;
        RECT 3.090 2.565 3.580 2.735 ;
        RECT 2.370 2.025 2.805 2.355 ;
        RECT 2.975 1.855 3.240 2.355 ;
        RECT 1.955 1.685 3.240 1.855 ;
        RECT 2.975 1.455 3.240 1.685 ;
        RECT 3.410 1.795 3.580 2.565 ;
        RECT 3.750 2.135 4.000 2.735 ;
        RECT 4.200 2.490 4.530 2.905 ;
        RECT 5.040 2.660 5.370 3.245 ;
        RECT 5.570 2.490 5.820 2.980 ;
        RECT 6.020 2.660 6.350 3.245 ;
        RECT 4.200 2.320 6.450 2.490 ;
        RECT 4.200 2.305 4.815 2.320 ;
        RECT 3.750 1.965 4.475 2.135 ;
        RECT 3.410 1.625 4.135 1.795 ;
        RECT 2.975 1.125 3.465 1.455 ;
        RECT 3.635 1.395 4.135 1.625 ;
        RECT 1.585 0.840 2.750 1.010 ;
        RECT 3.635 0.955 3.805 1.395 ;
        RECT 4.305 1.165 4.475 1.965 ;
        RECT 1.585 0.575 1.865 0.840 ;
        RECT 2.045 0.085 2.410 0.670 ;
        RECT 2.580 0.425 2.750 0.840 ;
        RECT 2.950 0.785 3.805 0.955 ;
        RECT 3.975 0.995 4.475 1.165 ;
        RECT 4.645 1.165 4.815 2.305 ;
        RECT 5.435 1.960 5.635 2.150 ;
        RECT 5.435 1.675 5.850 1.960 ;
        RECT 6.120 1.675 6.450 2.320 ;
        RECT 6.860 2.100 7.415 2.980 ;
        RECT 7.905 2.970 8.270 3.245 ;
        RECT 8.500 2.800 8.830 2.980 ;
        RECT 9.035 2.970 9.365 3.245 ;
        RECT 9.990 2.800 10.320 2.980 ;
        RECT 4.985 1.505 5.265 1.665 ;
        RECT 6.710 1.560 7.075 1.930 ;
        RECT 7.245 1.900 7.415 2.100 ;
        RECT 7.890 2.630 10.320 2.800 ;
        RECT 11.045 2.630 11.375 3.245 ;
        RECT 7.890 2.070 8.220 2.630 ;
        RECT 9.990 2.460 10.320 2.630 ;
        RECT 8.390 2.290 9.400 2.460 ;
        RECT 9.990 2.290 11.385 2.460 ;
        RECT 8.390 1.900 8.560 2.290 ;
        RECT 9.230 2.120 9.400 2.290 ;
        RECT 7.245 1.730 8.560 1.900 ;
        RECT 4.985 1.335 6.485 1.505 ;
        RECT 4.645 0.995 5.145 1.165 ;
        RECT 2.950 0.595 3.280 0.785 ;
        RECT 3.975 0.615 4.145 0.995 ;
        RECT 3.460 0.425 4.145 0.615 ;
        RECT 2.580 0.255 4.145 0.425 ;
        RECT 4.315 0.425 4.645 0.825 ;
        RECT 4.815 0.715 5.145 0.995 ;
        RECT 5.315 0.425 5.645 1.035 ;
        RECT 4.315 0.255 5.645 0.425 ;
        RECT 5.815 0.085 6.145 1.035 ;
        RECT 6.315 0.510 6.485 1.335 ;
        RECT 6.710 1.180 7.865 1.560 ;
        RECT 8.035 1.010 8.205 1.730 ;
        RECT 8.730 1.275 9.060 2.120 ;
        RECT 9.230 1.950 10.170 2.120 ;
        RECT 9.300 1.105 9.630 1.560 ;
        RECT 9.840 1.420 10.170 1.950 ;
        RECT 10.345 1.950 10.850 2.120 ;
        RECT 10.345 1.105 10.515 1.950 ;
        RECT 11.215 1.650 11.385 2.290 ;
        RECT 11.215 1.320 11.585 1.650 ;
        RECT 12.110 1.585 12.360 2.910 ;
        RECT 12.555 1.820 12.805 3.245 ;
        RECT 6.720 0.680 8.205 1.010 ;
        RECT 8.375 0.935 10.890 1.105 ;
        RECT 8.375 0.510 8.545 0.935 ;
        RECT 11.215 0.765 11.385 1.320 ;
        RECT 6.315 0.340 8.545 0.510 ;
        RECT 8.715 0.085 8.885 0.765 ;
        RECT 9.065 0.425 9.315 0.765 ;
        RECT 9.495 0.595 11.385 0.765 ;
        RECT 12.110 1.255 12.835 1.585 ;
        RECT 9.065 0.255 10.360 0.425 ;
        RECT 11.055 0.085 11.385 0.425 ;
        RECT 12.110 0.350 12.360 1.255 ;
        RECT 12.580 0.085 12.830 0.810 ;
        RECT 0.000 -0.085 13.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 3.035 1.210 3.205 1.380 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 8.795 1.950 8.965 2.120 ;
        RECT 6.875 1.210 7.045 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
      LAYER met1 ;
        RECT 2.975 1.365 3.265 1.410 ;
        RECT 6.815 1.365 7.105 1.410 ;
        RECT 2.975 1.225 7.105 1.365 ;
        RECT 2.975 1.180 3.265 1.225 ;
        RECT 6.815 1.180 7.105 1.225 ;
  END
END sky130_fd_sc_hs__dfbbn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfbbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.495 1.780 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.955 1.180 2.755 1.510 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 10.715 1.350 11.115 1.780 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER met1 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 8.735 2.105 9.025 2.150 ;
        RECT 5.375 1.965 9.025 2.105 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 8.735 1.920 9.025 1.965 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.205 1.240 6.580 1.305 ;
        RECT 10.555 1.240 12.515 1.370 ;
        RECT 0.005 1.145 1.415 1.240 ;
        RECT 4.205 1.145 14.395 1.240 ;
        RECT 0.005 0.245 14.395 1.145 ;
        RECT 0.000 0.000 14.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.400 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 13.515 1.940 13.845 2.980 ;
        RECT 13.515 1.770 14.035 1.940 ;
        RECT 13.865 1.100 14.035 1.770 ;
        RECT 13.540 0.850 14.035 1.100 ;
        RECT 13.540 0.350 13.800 0.850 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 11.645 2.020 11.815 2.980 ;
        RECT 11.645 1.850 11.985 2.020 ;
        RECT 11.815 1.180 11.985 1.850 ;
        RECT 11.630 0.440 11.985 1.180 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.400 3.415 ;
        RECT 0.105 2.120 0.435 2.980 ;
        RECT 0.635 2.290 0.805 3.245 ;
        RECT 1.005 2.905 2.125 3.075 ;
        RECT 0.105 1.950 0.835 2.120 ;
        RECT 0.665 1.630 0.835 1.950 ;
        RECT 1.005 1.820 1.445 2.905 ;
        RECT 0.665 1.300 1.105 1.630 ;
        RECT 0.665 1.130 0.835 1.300 ;
        RECT 1.275 1.130 1.445 1.820 ;
        RECT 0.115 0.960 0.835 1.130 ;
        RECT 0.115 0.350 0.365 0.960 ;
        RECT 0.545 0.085 0.875 0.790 ;
        RECT 1.055 0.350 1.445 1.130 ;
        RECT 1.615 1.010 1.785 2.735 ;
        RECT 1.955 1.855 2.125 2.905 ;
        RECT 2.295 2.525 2.465 3.245 ;
        RECT 2.635 2.905 4.605 3.075 ;
        RECT 2.635 2.355 2.805 2.905 ;
        RECT 3.085 2.565 3.570 2.735 ;
        RECT 2.365 2.025 2.805 2.355 ;
        RECT 2.975 1.855 3.230 2.355 ;
        RECT 1.955 1.685 3.230 1.855 ;
        RECT 3.005 1.455 3.230 1.685 ;
        RECT 3.400 1.795 3.570 2.565 ;
        RECT 3.740 2.135 3.990 2.735 ;
        RECT 4.185 2.490 4.605 2.905 ;
        RECT 5.055 2.660 5.385 3.245 ;
        RECT 5.565 2.490 5.895 2.980 ;
        RECT 6.095 2.660 6.425 3.245 ;
        RECT 4.185 2.320 6.380 2.490 ;
        RECT 4.185 2.305 4.775 2.320 ;
        RECT 3.740 1.965 4.435 2.135 ;
        RECT 3.400 1.625 4.095 1.795 ;
        RECT 3.715 1.465 4.095 1.625 ;
        RECT 3.005 1.125 3.545 1.455 ;
        RECT 1.615 0.840 2.780 1.010 ;
        RECT 3.715 0.955 3.885 1.465 ;
        RECT 4.265 1.295 4.435 1.965 ;
        RECT 1.615 0.575 1.865 0.840 ;
        RECT 2.045 0.085 2.440 0.670 ;
        RECT 2.610 0.425 2.780 0.840 ;
        RECT 2.980 0.785 3.885 0.955 ;
        RECT 4.055 1.125 4.435 1.295 ;
        RECT 4.605 1.295 4.775 2.305 ;
        RECT 4.945 1.610 5.245 1.940 ;
        RECT 5.415 1.630 5.745 2.150 ;
        RECT 6.050 1.630 6.380 2.320 ;
        RECT 6.965 2.100 7.455 2.980 ;
        RECT 8.010 2.970 8.340 3.245 ;
        RECT 8.570 2.800 8.900 2.980 ;
        RECT 9.105 2.970 9.435 3.245 ;
        RECT 10.060 2.800 10.390 2.980 ;
        RECT 5.075 1.460 5.245 1.610 ;
        RECT 4.605 1.125 4.905 1.295 ;
        RECT 5.075 1.290 6.415 1.460 ;
        RECT 2.980 0.595 3.310 0.785 ;
        RECT 4.055 0.615 4.225 1.125 ;
        RECT 4.735 1.120 4.905 1.125 ;
        RECT 3.490 0.425 4.225 0.615 ;
        RECT 2.610 0.255 4.225 0.425 ;
        RECT 4.395 0.435 4.565 0.955 ;
        RECT 4.735 0.605 5.075 1.120 ;
        RECT 5.245 0.435 5.575 1.025 ;
        RECT 4.395 0.265 5.575 0.435 ;
        RECT 5.745 0.085 6.075 1.025 ;
        RECT 6.245 0.510 6.415 1.290 ;
        RECT 6.785 1.410 7.115 1.910 ;
        RECT 7.285 1.890 7.455 2.100 ;
        RECT 7.925 2.630 10.390 2.800 ;
        RECT 11.115 2.630 11.445 3.245 ;
        RECT 7.925 2.060 8.255 2.630 ;
        RECT 10.060 2.460 10.390 2.630 ;
        RECT 8.425 2.290 9.890 2.460 ;
        RECT 10.060 2.290 11.460 2.460 ;
        RECT 8.425 1.890 8.595 2.290 ;
        RECT 7.285 1.720 8.595 1.890 ;
        RECT 8.765 1.780 8.995 2.120 ;
        RECT 9.720 1.890 9.890 2.290 ;
        RECT 10.375 1.950 10.920 2.120 ;
        RECT 7.685 1.410 7.935 1.550 ;
        RECT 6.785 1.180 7.935 1.410 ;
        RECT 8.105 1.010 8.275 1.720 ;
        RECT 8.765 1.450 9.160 1.780 ;
        RECT 9.720 1.720 10.205 1.890 ;
        RECT 9.370 1.180 9.700 1.550 ;
        RECT 9.910 1.470 10.205 1.720 ;
        RECT 10.375 1.180 10.545 1.950 ;
        RECT 11.290 1.680 11.460 2.290 ;
        RECT 12.015 2.190 12.345 3.245 ;
        RECT 12.545 1.820 12.875 2.860 ;
        RECT 13.065 1.820 13.315 3.245 ;
        RECT 14.045 2.110 14.295 3.245 ;
        RECT 11.290 1.350 11.645 1.680 ;
        RECT 12.635 1.600 12.875 1.820 ;
        RECT 6.650 0.680 8.275 1.010 ;
        RECT 8.445 1.010 10.990 1.180 ;
        RECT 8.445 0.510 8.615 1.010 ;
        RECT 11.290 0.840 11.460 1.350 ;
        RECT 12.635 1.270 13.695 1.600 ;
        RECT 6.245 0.340 8.615 0.510 ;
        RECT 8.785 0.085 8.955 0.840 ;
        RECT 9.135 0.425 9.385 0.840 ;
        RECT 9.605 0.670 11.460 0.840 ;
        RECT 9.605 0.595 9.935 0.670 ;
        RECT 10.110 0.425 10.440 0.500 ;
        RECT 9.135 0.255 10.440 0.425 ;
        RECT 10.665 0.085 11.450 0.500 ;
        RECT 12.155 0.085 12.405 1.260 ;
        RECT 12.635 0.350 12.885 1.270 ;
        RECT 13.095 0.085 13.370 1.050 ;
        RECT 13.970 0.085 14.300 0.680 ;
        RECT 0.000 -0.085 14.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 3.035 1.210 3.205 1.380 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 8.795 1.950 8.965 2.120 ;
        RECT 6.875 1.210 7.045 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
      LAYER met1 ;
        RECT 2.975 1.365 3.265 1.410 ;
        RECT 6.815 1.365 7.105 1.410 ;
        RECT 2.975 1.225 7.105 1.365 ;
        RECT 2.975 1.180 3.265 1.225 ;
        RECT 6.815 1.180 7.105 1.225 ;
  END
END sky130_fd_sc_hs__dfbbn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfbbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.180 0.805 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.960 1.825 2.290 2.155 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 10.235 0.980 10.580 1.650 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER li1 ;
        RECT 4.360 2.905 5.330 3.075 ;
        RECT 4.360 1.655 4.530 2.905 ;
        RECT 5.160 2.335 5.330 2.905 ;
        RECT 6.040 2.905 7.450 3.075 ;
        RECT 6.040 2.335 6.210 2.905 ;
        RECT 5.160 2.165 6.210 2.335 ;
        RECT 7.280 1.910 7.450 2.905 ;
        RECT 7.280 1.800 8.515 1.910 ;
        RECT 7.280 1.740 8.570 1.800 ;
        RECT 4.230 1.410 4.560 1.655 ;
        RECT 8.240 1.470 8.570 1.740 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.830 1.240 7.360 1.275 ;
        RECT 0.005 1.175 1.485 1.240 ;
        RECT 0.005 1.145 2.505 1.175 ;
        RECT 3.830 1.145 12.955 1.240 ;
        RECT 0.005 0.245 12.955 1.145 ;
        RECT 0.000 0.000 12.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.150 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.960 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.519000 ;
    PORT
      LAYER li1 ;
        RECT 12.525 0.350 12.860 2.980 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518900 ;
    PORT
      LAYER li1 ;
        RECT 11.120 1.820 11.460 2.980 ;
        RECT 11.290 1.130 11.460 1.820 ;
        RECT 11.065 0.350 11.460 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.085 1.890 0.535 2.980 ;
        RECT 0.705 2.060 1.035 3.245 ;
        RECT 0.085 1.720 1.145 1.890 ;
        RECT 0.085 1.010 0.255 1.720 ;
        RECT 0.975 1.300 1.145 1.720 ;
        RECT 1.315 1.585 1.565 2.980 ;
        RECT 1.805 2.425 2.410 3.245 ;
        RECT 2.580 2.295 2.955 2.755 ;
        RECT 1.315 1.255 2.615 1.585 ;
        RECT 1.315 1.130 1.485 1.255 ;
        RECT 0.085 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 1.010 ;
        RECT 1.125 0.350 1.485 1.130 ;
        RECT 2.785 1.085 2.955 2.295 ;
        RECT 1.655 0.085 1.905 1.065 ;
        RECT 2.085 0.915 2.955 1.085 ;
        RECT 3.125 1.795 3.430 2.335 ;
        RECT 3.940 1.965 4.190 3.245 ;
        RECT 4.700 1.995 4.950 2.735 ;
        RECT 5.500 2.505 5.870 3.245 ;
        RECT 6.540 2.280 6.870 2.735 ;
        RECT 7.620 2.650 8.420 3.245 ;
        RECT 8.685 2.410 8.935 2.980 ;
        RECT 9.470 2.580 9.800 3.245 ;
        RECT 10.590 2.580 10.920 3.245 ;
        RECT 8.685 2.380 10.950 2.410 ;
        RECT 6.540 2.110 7.110 2.280 ;
        RECT 4.700 1.825 6.020 1.995 ;
        RECT 3.125 1.625 4.060 1.795 ;
        RECT 2.085 0.605 2.335 0.915 ;
        RECT 3.125 0.745 3.295 1.625 ;
        RECT 2.575 0.415 3.295 0.745 ;
        RECT 3.465 0.900 3.720 1.455 ;
        RECT 3.890 1.240 4.060 1.625 ;
        RECT 5.850 1.585 6.020 1.825 ;
        RECT 6.440 1.610 6.770 1.940 ;
        RECT 4.745 1.255 5.100 1.585 ;
        RECT 4.745 1.240 4.915 1.255 ;
        RECT 3.890 1.070 4.915 1.240 ;
        RECT 5.310 1.180 5.640 1.585 ;
        RECT 5.850 1.255 6.180 1.585 ;
        RECT 5.850 1.010 6.020 1.255 ;
        RECT 5.085 0.900 6.020 1.010 ;
        RECT 3.465 0.840 6.020 0.900 ;
        RECT 3.465 0.730 5.335 0.840 ;
        RECT 5.015 0.595 5.335 0.730 ;
        RECT 6.190 0.670 6.430 1.085 ;
        RECT 3.560 0.085 4.155 0.560 ;
        RECT 4.415 0.425 4.825 0.560 ;
        RECT 5.510 0.425 5.840 0.670 ;
        RECT 4.415 0.255 5.840 0.425 ;
        RECT 6.060 0.085 6.430 0.670 ;
        RECT 6.600 0.425 6.770 1.610 ;
        RECT 6.940 1.570 7.110 2.110 ;
        RECT 7.620 2.240 10.950 2.380 ;
        RECT 7.620 2.080 9.385 2.240 ;
        RECT 8.685 1.970 9.385 2.080 ;
        RECT 6.940 1.400 8.070 1.570 ;
        RECT 6.940 0.595 7.175 1.400 ;
        RECT 7.900 1.300 8.070 1.400 ;
        RECT 8.780 1.300 9.045 1.550 ;
        RECT 7.345 0.425 7.670 1.230 ;
        RECT 7.900 1.130 9.045 1.300 ;
        RECT 9.215 0.960 9.385 1.970 ;
        RECT 9.710 1.820 10.405 2.070 ;
        RECT 9.710 1.190 10.065 1.820 ;
        RECT 10.780 1.650 10.950 2.240 ;
        RECT 11.640 2.030 11.890 2.910 ;
        RECT 10.780 1.320 11.120 1.650 ;
        RECT 11.640 1.585 11.810 2.030 ;
        RECT 12.075 1.820 12.325 3.245 ;
        RECT 6.600 0.255 7.670 0.425 ;
        RECT 8.085 0.085 8.415 0.960 ;
        RECT 8.585 0.425 8.915 0.960 ;
        RECT 9.085 0.595 9.385 0.960 ;
        RECT 9.555 0.425 9.725 1.020 ;
        RECT 8.585 0.255 9.725 0.425 ;
        RECT 9.895 0.810 10.065 1.190 ;
        RECT 11.640 1.255 12.355 1.585 ;
        RECT 9.895 0.350 10.385 0.810 ;
        RECT 10.565 0.085 10.895 0.810 ;
        RECT 11.640 0.350 11.875 1.255 ;
        RECT 12.055 0.085 12.305 0.810 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 5.435 1.210 5.605 1.380 ;
        RECT 9.755 1.210 9.925 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
      LAYER met1 ;
        RECT 5.375 1.365 5.665 1.410 ;
        RECT 9.695 1.365 9.985 1.410 ;
        RECT 5.375 1.225 9.985 1.365 ;
        RECT 5.375 1.180 5.665 1.225 ;
        RECT 9.695 1.180 9.985 1.225 ;
  END
END sky130_fd_sc_hs__dfbbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.640 2.275 1.780 ;
        RECT 1.810 1.310 2.275 1.640 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.000 0.520 2.195 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 2.105 1.345 2.150 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 1.055 1.965 8.065 2.105 ;
        RECT 1.055 1.920 1.345 1.965 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.520 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.480 1.140 3.030 1.240 ;
        RECT 5.475 1.140 6.025 1.280 ;
        RECT 1.480 0.940 6.500 1.140 ;
        RECT 0.060 0.920 6.500 0.940 ;
        RECT 8.950 0.920 11.505 1.240 ;
        RECT 0.060 0.245 11.505 0.920 ;
        RECT 0.000 0.000 11.520 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.710 3.520 ;
        RECT 1.415 1.620 7.060 1.660 ;
        RECT 5.540 1.555 7.060 1.620 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.520 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 11.075 1.820 11.435 2.980 ;
        RECT 11.265 1.130 11.435 1.820 ;
        RECT 11.065 0.350 11.435 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.951500 ;
    PORT
      LAYER li1 ;
        RECT 9.260 1.810 9.950 2.985 ;
        RECT 9.560 0.350 9.950 1.810 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.115 2.520 0.365 3.245 ;
        RECT 0.565 2.520 0.895 2.980 ;
        RECT 1.095 2.650 1.345 3.245 ;
        RECT 2.025 2.650 2.355 3.245 ;
        RECT 4.440 2.755 4.785 3.245 ;
        RECT 0.690 2.480 0.895 2.520 ;
        RECT 3.065 2.480 3.395 2.755 ;
        RECT 0.690 2.310 3.395 2.480 ;
        RECT 3.595 2.585 3.845 2.755 ;
        RECT 4.990 2.585 5.325 2.680 ;
        RECT 3.595 2.415 5.325 2.585 ;
        RECT 0.690 0.830 0.860 2.310 ;
        RECT 3.065 2.245 3.395 2.310 ;
        RECT 1.030 1.130 1.300 2.140 ;
        RECT 1.470 1.810 1.825 2.140 ;
        RECT 2.475 1.905 2.805 2.140 ;
        RECT 3.065 2.075 3.840 2.245 ;
        RECT 1.470 1.140 1.640 1.810 ;
        RECT 2.475 1.735 3.500 1.905 ;
        RECT 2.945 1.575 3.500 1.735 ;
        RECT 2.445 1.140 2.775 1.550 ;
        RECT 1.470 0.970 2.775 1.140 ;
        RECT 0.170 0.660 0.860 0.830 ;
        RECT 0.170 0.370 0.500 0.660 ;
        RECT 1.030 0.085 1.280 0.830 ;
        RECT 1.470 0.350 1.920 0.970 ;
        RECT 2.945 0.800 3.115 1.575 ;
        RECT 3.670 1.370 3.840 2.075 ;
        RECT 2.090 0.085 2.420 0.800 ;
        RECT 2.590 0.425 3.115 0.800 ;
        RECT 3.285 1.200 3.840 1.370 ;
        RECT 3.285 0.595 3.535 1.200 ;
        RECT 4.010 1.030 4.180 2.415 ;
        RECT 4.890 2.350 5.325 2.415 ;
        RECT 3.705 0.595 4.180 1.030 ;
        RECT 4.350 1.090 4.630 2.155 ;
        RECT 4.890 1.615 5.060 2.350 ;
        RECT 5.230 1.825 5.610 2.155 ;
        RECT 5.780 1.740 6.030 3.245 ;
        RECT 4.890 1.445 5.560 1.615 ;
        RECT 6.230 1.570 6.480 2.755 ;
        RECT 6.700 2.365 7.665 2.695 ;
        RECT 5.230 1.285 5.560 1.445 ;
        RECT 5.745 1.400 6.480 1.570 ;
        RECT 6.650 1.865 7.325 2.195 ;
        RECT 5.745 1.090 5.915 1.400 ;
        RECT 6.650 1.230 6.820 1.865 ;
        RECT 7.495 1.595 7.665 2.365 ;
        RECT 7.835 2.335 8.060 3.245 ;
        RECT 8.260 2.335 8.640 2.730 ;
        RECT 7.835 1.835 8.300 2.165 ;
        RECT 8.470 1.935 8.640 2.335 ;
        RECT 8.810 2.105 9.025 3.245 ;
        RECT 8.470 1.765 8.970 1.935 ;
        RECT 4.350 0.920 5.915 1.090 ;
        RECT 6.085 0.900 6.820 1.230 ;
        RECT 6.990 1.425 8.630 1.595 ;
        RECT 6.085 0.750 6.255 0.900 ;
        RECT 4.350 0.580 6.255 0.750 ;
        RECT 6.990 0.730 7.160 1.425 ;
        RECT 8.330 1.265 8.630 1.425 ;
        RECT 7.430 1.070 7.760 1.230 ;
        RECT 8.800 1.070 8.970 1.765 ;
        RECT 10.190 1.630 10.440 2.975 ;
        RECT 10.610 1.820 10.905 3.245 ;
        RECT 10.190 1.300 11.095 1.630 ;
        RECT 7.430 0.900 8.970 1.070 ;
        RECT 4.350 0.425 4.520 0.580 ;
        RECT 2.590 0.255 4.520 0.425 ;
        RECT 4.995 0.085 5.325 0.410 ;
        RECT 6.425 0.400 7.160 0.730 ;
        RECT 7.535 0.085 7.995 0.680 ;
        RECT 8.485 0.350 8.970 0.900 ;
        RECT 9.140 0.085 9.390 1.130 ;
        RECT 10.190 0.350 10.440 1.300 ;
        RECT 10.645 0.085 10.895 1.130 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
  END
END sky130_fd_sc_hs__dfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 6.705 1.180 7.045 1.670 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.810 0.515 1.570 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.735 1.345 1.780 ;
        RECT 2.495 1.735 2.785 1.780 ;
        RECT 9.695 1.735 9.985 1.780 ;
        RECT 1.055 1.595 9.985 1.735 ;
        RECT 1.055 1.550 1.345 1.595 ;
        RECT 2.495 1.550 2.785 1.595 ;
        RECT 9.695 1.550 9.985 1.595 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.380 1.570 4.990 1.710 ;
        RECT 3.235 1.360 4.990 1.570 ;
        RECT 3.235 1.295 7.070 1.360 ;
        RECT 1.140 0.955 2.085 1.240 ;
        RECT 3.235 0.955 8.875 1.295 ;
        RECT 1.140 0.920 8.875 0.955 ;
        RECT 10.655 0.920 13.915 1.240 ;
        RECT 0.220 0.245 13.915 0.920 ;
        RECT 0.000 0.000 13.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 2.245 14.110 3.520 ;
        RECT -0.190 1.660 3.025 2.245 ;
        RECT 5.200 1.660 14.110 2.245 ;
        RECT 10.235 1.580 12.385 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.920 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 12.975 1.820 13.305 2.980 ;
        RECT 13.135 1.130 13.305 1.820 ;
        RECT 13.060 0.330 13.390 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 10.895 1.540 11.065 2.900 ;
        RECT 10.895 1.410 11.725 1.540 ;
        RECT 10.895 1.320 11.875 1.410 ;
        RECT 11.195 0.770 11.875 1.320 ;
        RECT 11.195 0.350 11.455 0.770 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.920 3.415 ;
        RECT 0.115 2.965 1.435 3.245 ;
        RECT 0.115 1.940 0.510 2.965 ;
        RECT 1.605 2.905 2.775 3.075 ;
        RECT 1.605 2.795 1.775 2.905 ;
        RECT 0.680 2.625 1.775 2.795 ;
        RECT 0.680 1.950 1.010 2.625 ;
        RECT 1.485 2.285 1.970 2.455 ;
        RECT 0.685 0.640 0.855 1.950 ;
        RECT 1.025 1.450 1.315 1.780 ;
        RECT 1.485 1.185 1.655 2.285 ;
        RECT 2.185 2.115 2.435 2.735 ;
        RECT 2.605 2.455 2.775 2.905 ;
        RECT 2.945 2.625 3.195 3.245 ;
        RECT 3.365 2.905 4.460 3.075 ;
        RECT 3.365 2.455 3.535 2.905 ;
        RECT 4.290 2.815 4.460 2.905 ;
        RECT 2.605 2.285 3.535 2.455 ;
        RECT 3.790 2.115 4.120 2.735 ;
        RECT 4.290 2.485 4.960 2.815 ;
        RECT 5.425 2.595 5.785 2.980 ;
        RECT 5.990 2.765 6.500 3.245 ;
        RECT 7.315 2.905 8.220 3.075 ;
        RECT 7.315 2.595 7.505 2.905 ;
        RECT 4.290 2.410 4.475 2.485 ;
        RECT 1.825 1.945 4.120 2.115 ;
        RECT 1.825 1.470 2.155 1.945 ;
        RECT 2.385 1.445 2.755 1.775 ;
        RECT 2.925 1.555 3.255 1.775 ;
        RECT 3.885 1.610 4.120 1.945 ;
        RECT 2.925 1.185 3.095 1.555 ;
        RECT 1.485 1.015 3.095 1.185 ;
        RECT 3.345 1.105 3.715 1.385 ;
        RECT 3.885 1.275 4.135 1.610 ;
        RECT 4.305 1.105 4.475 2.410 ;
        RECT 5.425 2.425 7.505 2.595 ;
        RECT 5.425 2.240 5.785 2.425 ;
        RECT 4.645 1.910 5.785 2.240 ;
        RECT 6.705 2.170 7.035 2.255 ;
        RECT 5.095 1.840 5.785 1.910 ;
        RECT 6.095 1.840 7.505 2.170 ;
        RECT 0.325 0.390 0.855 0.640 ;
        RECT 1.145 0.085 1.475 0.810 ;
        RECT 1.645 0.350 1.975 1.015 ;
        RECT 2.205 0.085 2.535 0.780 ;
        RECT 2.705 0.425 2.875 1.015 ;
        RECT 3.345 0.935 4.475 1.105 ;
        RECT 4.645 0.765 4.895 1.600 ;
        RECT 5.095 1.000 5.425 1.840 ;
        RECT 6.095 1.670 6.265 1.840 ;
        RECT 5.595 1.340 6.535 1.670 ;
        RECT 7.710 1.525 7.880 2.735 ;
        RECT 6.365 0.965 6.535 1.340 ;
        RECT 7.215 1.355 7.880 1.525 ;
        RECT 8.050 1.605 8.220 2.905 ;
        RECT 8.390 2.095 8.640 2.385 ;
        RECT 9.265 2.290 9.625 3.245 ;
        RECT 9.830 2.120 10.160 2.385 ;
        RECT 10.365 2.290 10.695 3.245 ;
        RECT 8.390 1.925 8.895 2.095 ;
        RECT 3.045 0.595 4.895 0.765 ;
        RECT 5.065 0.660 6.195 0.830 ;
        RECT 5.065 0.425 5.235 0.660 ;
        RECT 2.705 0.255 5.235 0.425 ;
        RECT 5.605 0.085 5.855 0.490 ;
        RECT 6.025 0.425 6.195 0.660 ;
        RECT 6.365 0.635 6.960 0.965 ;
        RECT 7.215 0.425 7.385 1.355 ;
        RECT 8.050 1.275 8.555 1.605 ;
        RECT 8.725 1.265 8.895 1.925 ;
        RECT 9.065 1.950 10.675 2.120 ;
        RECT 9.065 1.455 9.330 1.950 ;
        RECT 9.540 1.450 9.955 1.780 ;
        RECT 7.555 0.765 7.725 1.185 ;
        RECT 8.725 1.105 10.335 1.265 ;
        RECT 7.905 0.935 10.335 1.105 ;
        RECT 10.505 0.765 10.675 1.950 ;
        RECT 11.265 1.740 11.595 3.245 ;
        RECT 11.895 1.740 12.305 2.780 ;
        RECT 12.475 1.820 12.805 3.245 ;
        RECT 13.475 1.820 13.805 3.245 ;
        RECT 12.135 1.630 12.305 1.740 ;
        RECT 12.135 1.300 12.965 1.630 ;
        RECT 7.555 0.595 9.235 0.765 ;
        RECT 6.025 0.255 8.780 0.425 ;
        RECT 8.985 0.350 9.235 0.595 ;
        RECT 9.415 0.085 9.745 0.720 ;
        RECT 10.205 0.350 10.675 0.765 ;
        RECT 10.845 0.085 11.015 1.100 ;
        RECT 11.625 0.085 11.965 0.600 ;
        RECT 12.135 0.350 12.430 1.300 ;
        RECT 12.630 0.085 12.880 1.130 ;
        RECT 13.560 0.085 13.820 1.130 ;
        RECT 0.000 -0.085 13.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 1.115 1.580 1.285 1.750 ;
        RECT 2.555 1.580 2.725 1.750 ;
        RECT 9.755 1.580 9.925 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
  END
END sky130_fd_sc_hs__dfrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.180 1.765 1.550 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.960 0.370 2.150 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.735 1.345 1.780 ;
        RECT 4.895 1.735 5.185 1.780 ;
        RECT 8.255 1.735 8.545 1.780 ;
        RECT 1.055 1.595 8.545 1.735 ;
        RECT 1.055 1.550 1.345 1.595 ;
        RECT 4.895 1.550 5.185 1.595 ;
        RECT 8.255 1.550 8.545 1.595 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.495 1.370 3.015 1.415 ;
        RECT 1.915 1.240 3.015 1.370 ;
        RECT 0.935 1.185 3.015 1.240 ;
        RECT 5.360 1.185 6.710 1.465 ;
        RECT 0.935 1.145 6.710 1.185 ;
        RECT 10.050 1.150 11.035 1.340 ;
        RECT 9.540 1.145 11.035 1.150 ;
        RECT 0.935 0.920 11.035 1.145 ;
        RECT 0.035 0.245 11.035 0.920 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.675 11.230 3.520 ;
        RECT -0.190 1.660 3.225 1.675 ;
        RECT 6.920 1.660 11.230 1.675 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.533800 ;
    PORT
      LAYER li1 ;
        RECT 10.605 1.820 10.955 2.980 ;
        RECT 10.785 1.150 10.955 1.820 ;
        RECT 10.590 0.440 10.955 1.150 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.110 2.520 0.440 3.245 ;
        RECT 0.640 2.350 0.890 2.980 ;
        RECT 1.060 2.655 1.390 3.245 ;
        RECT 2.070 2.655 2.400 3.245 ;
        RECT 3.170 2.485 3.420 2.980 ;
        RECT 3.620 2.520 4.055 2.980 ;
        RECT 4.460 2.520 4.790 3.245 ;
        RECT 1.060 2.350 3.420 2.485 ;
        RECT 0.540 2.315 3.420 2.350 ;
        RECT 0.540 2.180 1.230 2.315 ;
        RECT 0.540 0.790 0.710 2.180 ;
        RECT 1.515 1.820 2.165 2.145 ;
        RECT 0.880 1.350 1.285 1.780 ;
        RECT 1.935 1.010 2.165 1.820 ;
        RECT 0.145 0.350 0.710 0.790 ;
        RECT 1.045 0.085 1.295 0.810 ;
        RECT 1.475 0.635 2.165 1.010 ;
        RECT 2.335 0.805 2.505 2.315 ;
        RECT 3.885 2.190 4.055 2.520 ;
        RECT 4.970 2.190 5.300 2.980 ;
        RECT 5.490 2.360 5.820 3.245 ;
        RECT 2.675 2.105 2.940 2.145 ;
        RECT 2.675 1.775 3.715 2.105 ;
        RECT 3.885 2.020 5.695 2.190 ;
        RECT 5.990 2.140 6.700 2.980 ;
        RECT 6.870 2.705 7.600 2.865 ;
        RECT 6.870 2.535 7.900 2.705 ;
        RECT 2.675 1.415 2.940 1.775 ;
        RECT 2.675 1.245 3.705 1.415 ;
        RECT 2.675 0.975 2.940 1.245 ;
        RECT 3.115 0.805 3.365 1.075 ;
        RECT 2.335 0.635 3.365 0.805 ;
        RECT 1.475 0.350 1.805 0.635 ;
        RECT 3.535 0.465 3.705 1.245 ;
        RECT 3.885 1.075 4.055 2.020 ;
        RECT 4.280 1.520 4.610 1.850 ;
        RECT 4.440 1.300 4.610 1.520 ;
        RECT 4.820 1.470 5.155 1.800 ;
        RECT 5.365 1.470 5.695 2.020 ;
        RECT 5.865 1.970 6.700 2.140 ;
        RECT 5.865 1.300 6.035 1.970 ;
        RECT 7.310 1.800 7.560 2.365 ;
        RECT 6.205 1.630 7.560 1.800 ;
        RECT 6.205 1.470 6.510 1.630 ;
        RECT 4.440 1.130 6.195 1.300 ;
        RECT 6.750 1.295 7.420 1.455 ;
        RECT 3.875 0.635 4.125 1.075 ;
        RECT 4.295 0.790 5.695 0.960 ;
        RECT 4.295 0.465 4.465 0.790 ;
        RECT 2.020 0.085 2.350 0.465 ;
        RECT 3.035 0.255 4.465 0.465 ;
        RECT 5.025 0.085 5.355 0.620 ;
        RECT 5.525 0.425 5.695 0.790 ;
        RECT 5.865 0.595 6.195 1.130 ;
        RECT 6.365 1.125 7.420 1.295 ;
        RECT 7.730 1.295 7.900 2.535 ;
        RECT 8.140 2.520 8.470 3.245 ;
        RECT 8.680 2.335 9.010 2.980 ;
        RECT 9.210 2.520 9.460 3.245 ;
        RECT 8.070 2.135 9.050 2.335 ;
        RECT 9.650 2.305 9.980 2.980 ;
        RECT 8.070 1.965 9.560 2.135 ;
        RECT 8.285 1.465 8.710 1.795 ;
        RECT 8.920 1.295 9.220 1.795 ;
        RECT 7.730 1.125 9.220 1.295 ;
        RECT 6.365 0.425 6.535 1.125 ;
        RECT 7.730 0.955 7.900 1.125 ;
        RECT 9.390 0.955 9.560 1.965 ;
        RECT 6.705 0.625 7.900 0.955 ;
        RECT 5.525 0.255 6.535 0.425 ;
        RECT 8.115 0.085 8.555 0.905 ;
        RECT 9.045 0.575 9.560 0.955 ;
        RECT 9.730 1.650 9.980 2.305 ;
        RECT 10.150 2.100 10.400 3.245 ;
        RECT 9.730 1.320 10.615 1.650 ;
        RECT 9.730 0.530 9.980 1.320 ;
        RECT 10.160 0.085 10.410 1.130 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 1.115 1.580 1.285 1.750 ;
        RECT 4.955 1.580 5.125 1.750 ;
        RECT 8.315 1.580 8.485 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__dfrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.640 2.275 1.780 ;
        RECT 1.795 1.310 2.275 1.640 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.000 0.515 2.170 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 2.105 1.345 2.150 ;
        RECT 4.895 2.105 5.185 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 1.055 1.965 8.065 2.105 ;
        RECT 1.055 1.920 1.345 1.965 ;
        RECT 4.895 1.920 5.185 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.400 0.955 6.710 1.240 ;
        RECT 10.055 1.050 11.035 1.240 ;
        RECT 9.065 0.955 11.035 1.050 ;
        RECT 1.400 0.940 11.035 0.955 ;
        RECT 0.020 0.245 11.035 0.940 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
        RECT 1.390 1.650 6.400 1.660 ;
        RECT 5.320 1.555 6.400 1.650 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.591700 ;
    PORT
      LAYER li1 ;
        RECT 9.725 1.885 10.425 2.980 ;
        RECT 10.165 1.130 10.425 1.885 ;
        RECT 10.165 0.350 10.495 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.105 2.520 0.355 3.245 ;
        RECT 0.555 2.520 0.885 2.980 ;
        RECT 1.085 2.650 1.335 3.245 ;
        RECT 1.985 2.680 2.315 3.245 ;
        RECT 4.385 2.740 4.715 3.245 ;
        RECT 0.685 2.480 0.885 2.520 ;
        RECT 3.010 2.510 3.260 2.725 ;
        RECT 1.505 2.480 3.260 2.510 ;
        RECT 0.685 2.340 3.260 2.480 ;
        RECT 3.460 2.570 3.790 2.725 ;
        RECT 3.460 2.400 5.250 2.570 ;
        RECT 0.685 2.310 1.675 2.340 ;
        RECT 0.685 0.830 0.855 2.310 ;
        RECT 3.010 2.230 3.260 2.340 ;
        RECT 1.025 1.130 1.285 2.140 ;
        RECT 1.455 1.810 1.865 2.140 ;
        RECT 2.515 1.890 2.765 2.170 ;
        RECT 3.010 2.060 3.755 2.230 ;
        RECT 1.455 1.140 1.625 1.810 ;
        RECT 2.515 1.720 3.415 1.890 ;
        RECT 2.865 1.560 3.415 1.720 ;
        RECT 2.445 1.140 2.695 1.550 ;
        RECT 1.455 0.970 2.695 1.140 ;
        RECT 0.130 0.660 0.855 0.830 ;
        RECT 0.130 0.370 0.460 0.660 ;
        RECT 1.030 0.085 1.280 0.830 ;
        RECT 1.455 0.350 1.840 0.970 ;
        RECT 2.865 0.800 3.035 1.560 ;
        RECT 3.585 1.390 3.755 2.060 ;
        RECT 2.010 0.085 2.340 0.800 ;
        RECT 2.510 0.500 3.035 0.800 ;
        RECT 3.205 1.220 3.755 1.390 ;
        RECT 3.205 0.670 3.455 1.220 ;
        RECT 3.925 1.050 4.095 2.400 ;
        RECT 4.615 2.320 5.250 2.400 ;
        RECT 3.625 0.670 4.095 1.050 ;
        RECT 4.265 1.075 4.445 2.125 ;
        RECT 4.615 1.575 4.785 2.320 ;
        RECT 4.955 1.795 5.285 2.150 ;
        RECT 5.480 1.745 5.810 3.245 ;
        RECT 5.980 1.865 6.310 2.755 ;
        RECT 6.480 2.475 7.635 2.805 ;
        RECT 4.615 1.245 5.650 1.575 ;
        RECT 5.980 1.130 6.150 1.865 ;
        RECT 6.480 1.685 6.650 2.475 ;
        RECT 5.820 1.075 6.150 1.130 ;
        RECT 4.265 0.905 6.150 1.075 ;
        RECT 4.265 0.565 5.650 0.735 ;
        RECT 5.820 0.665 6.150 0.905 ;
        RECT 6.320 1.515 6.650 1.685 ;
        RECT 6.320 0.845 6.490 1.515 ;
        RECT 6.965 1.345 7.295 2.305 ;
        RECT 7.465 1.685 7.635 2.475 ;
        RECT 7.805 2.445 8.135 3.245 ;
        RECT 8.320 2.445 8.685 2.905 ;
        RECT 7.805 1.920 8.345 2.255 ;
        RECT 8.515 2.025 8.685 2.445 ;
        RECT 8.855 2.195 9.185 3.245 ;
        RECT 8.515 1.855 9.190 2.025 ;
        RECT 7.465 1.515 8.850 1.685 ;
        RECT 8.520 1.355 8.850 1.515 ;
        RECT 6.690 1.015 7.420 1.345 ;
        RECT 7.590 1.185 7.920 1.345 ;
        RECT 9.020 1.185 9.190 1.855 ;
        RECT 9.385 1.715 9.555 2.905 ;
        RECT 10.595 1.820 10.925 3.245 ;
        RECT 9.385 1.385 9.935 1.715 ;
        RECT 7.590 1.015 9.190 1.185 ;
        RECT 6.320 0.595 7.080 0.845 ;
        RECT 4.265 0.500 4.435 0.565 ;
        RECT 2.510 0.330 4.435 0.500 ;
        RECT 5.480 0.425 5.650 0.565 ;
        RECT 7.250 0.425 7.420 1.015 ;
        RECT 4.915 0.085 5.310 0.395 ;
        RECT 5.480 0.255 7.420 0.425 ;
        RECT 7.745 0.085 8.075 0.845 ;
        RECT 8.615 0.385 8.945 1.015 ;
        RECT 9.175 0.085 9.425 0.845 ;
        RECT 9.605 0.350 9.935 1.385 ;
        RECT 10.675 0.085 10.925 1.130 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 4.955 1.950 5.125 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__dfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.650 2.275 1.780 ;
        RECT 1.795 1.320 2.275 1.650 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.000 0.495 2.170 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 2.105 1.345 2.150 ;
        RECT 4.895 2.105 5.185 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 1.055 1.965 8.065 2.105 ;
        RECT 1.055 1.920 1.345 1.965 ;
        RECT 4.895 1.920 5.185 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.520 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.400 0.955 6.735 1.240 ;
        RECT 9.125 0.955 11.515 1.240 ;
        RECT 1.400 0.940 11.515 0.955 ;
        RECT 0.020 0.245 11.515 0.940 ;
        RECT 0.000 0.000 11.520 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.710 3.520 ;
        RECT 1.390 1.555 6.930 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.520 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 10.650 0.350 10.980 2.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.105 2.520 0.435 3.245 ;
        RECT 0.635 2.520 0.835 2.980 ;
        RECT 1.005 2.660 1.335 3.245 ;
        RECT 1.985 2.660 2.315 3.245 ;
        RECT 4.420 2.755 4.750 3.245 ;
        RECT 0.665 2.490 0.835 2.520 ;
        RECT 3.015 2.490 3.265 2.725 ;
        RECT 0.665 2.320 3.265 2.490 ;
        RECT 3.465 2.585 3.795 2.725 ;
        RECT 3.465 2.415 5.285 2.585 ;
        RECT 0.665 0.830 0.835 2.320 ;
        RECT 3.015 2.290 3.265 2.320 ;
        RECT 3.095 2.245 3.265 2.290 ;
        RECT 1.005 1.140 1.285 2.150 ;
        RECT 1.455 1.820 1.865 2.150 ;
        RECT 2.515 1.905 2.870 2.120 ;
        RECT 3.095 2.075 3.760 2.245 ;
        RECT 1.455 1.150 1.625 1.820 ;
        RECT 2.515 1.735 3.420 1.905 ;
        RECT 2.870 1.575 3.420 1.735 ;
        RECT 2.445 1.150 2.700 1.550 ;
        RECT 1.455 0.980 2.700 1.150 ;
        RECT 0.130 0.660 0.835 0.830 ;
        RECT 0.130 0.370 0.460 0.660 ;
        RECT 1.030 0.085 1.280 0.830 ;
        RECT 1.455 0.350 1.840 0.980 ;
        RECT 2.870 0.810 3.040 1.575 ;
        RECT 3.590 1.405 3.760 2.075 ;
        RECT 2.010 0.085 2.340 0.810 ;
        RECT 2.510 0.500 3.040 0.810 ;
        RECT 3.210 1.235 3.760 1.405 ;
        RECT 3.210 0.670 3.460 1.235 ;
        RECT 3.930 1.065 4.100 2.415 ;
        RECT 4.615 2.320 5.285 2.415 ;
        RECT 3.630 0.670 4.100 1.065 ;
        RECT 4.270 1.125 4.445 2.125 ;
        RECT 4.615 1.575 4.785 2.320 ;
        RECT 4.955 1.795 5.285 2.150 ;
        RECT 5.515 1.745 5.845 3.245 ;
        RECT 6.015 1.855 6.345 2.755 ;
        RECT 6.515 2.475 7.625 2.805 ;
        RECT 4.615 1.295 5.685 1.575 ;
        RECT 6.015 1.130 6.185 1.855 ;
        RECT 6.515 1.685 6.685 2.475 ;
        RECT 5.855 1.125 6.185 1.130 ;
        RECT 4.270 0.955 6.185 1.125 ;
        RECT 4.270 0.615 5.685 0.785 ;
        RECT 4.270 0.500 4.440 0.615 ;
        RECT 2.510 0.330 4.440 0.500 ;
        RECT 4.920 0.085 5.345 0.445 ;
        RECT 5.515 0.425 5.685 0.615 ;
        RECT 5.855 0.595 6.185 0.955 ;
        RECT 6.355 1.515 6.685 1.685 ;
        RECT 6.355 0.845 6.525 1.515 ;
        RECT 6.955 1.345 7.285 2.305 ;
        RECT 7.455 1.730 7.625 2.475 ;
        RECT 7.795 2.445 8.125 3.245 ;
        RECT 8.295 2.445 8.885 2.775 ;
        RECT 9.090 2.445 9.420 3.245 ;
        RECT 8.715 2.275 8.885 2.445 ;
        RECT 7.805 1.920 8.395 2.275 ;
        RECT 8.715 2.105 9.375 2.275 ;
        RECT 8.705 1.730 9.035 1.890 ;
        RECT 7.455 1.560 9.035 1.730 ;
        RECT 9.205 1.390 9.375 2.105 ;
        RECT 9.590 2.030 9.920 2.905 ;
        RECT 6.725 1.015 7.455 1.345 ;
        RECT 7.625 1.220 9.375 1.390 ;
        RECT 9.660 1.630 9.920 2.030 ;
        RECT 10.150 1.820 10.480 3.245 ;
        RECT 11.155 1.820 11.405 3.245 ;
        RECT 9.660 1.300 10.190 1.630 ;
        RECT 7.625 1.060 7.955 1.220 ;
        RECT 6.355 0.595 7.115 0.845 ;
        RECT 7.285 0.425 7.455 1.015 ;
        RECT 5.515 0.255 7.455 0.425 ;
        RECT 7.770 0.085 8.190 0.715 ;
        RECT 8.680 0.385 9.010 1.220 ;
        RECT 9.230 0.085 9.480 1.050 ;
        RECT 9.660 0.350 9.990 1.300 ;
        RECT 10.220 0.085 10.470 1.130 ;
        RECT 11.160 0.085 11.410 1.130 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 4.955 1.950 5.125 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
  END
END sky130_fd_sc_hs__dfrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.640 2.275 1.780 ;
        RECT 1.795 1.310 2.275 1.640 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.000 0.515 2.180 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 2.105 1.345 2.150 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 8.735 2.105 9.025 2.150 ;
        RECT 1.055 1.965 9.025 2.105 ;
        RECT 1.055 1.920 1.345 1.965 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 8.735 1.920 9.025 1.965 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.435 0.955 7.565 1.240 ;
        RECT 9.950 0.955 13.435 1.240 ;
        RECT 1.435 0.940 13.435 0.955 ;
        RECT 0.055 0.245 13.435 0.940 ;
        RECT 0.000 0.000 13.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.630 3.520 ;
        RECT 1.400 1.650 2.935 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.440 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.207100 ;
    PORT
      LAYER li1 ;
        RECT 11.035 1.970 11.365 2.980 ;
        RECT 12.410 1.970 12.740 2.980 ;
        RECT 11.035 1.800 12.740 1.970 ;
        RECT 12.410 1.780 12.740 1.800 ;
        RECT 12.410 1.610 13.315 1.780 ;
        RECT 12.575 1.270 13.315 1.610 ;
        RECT 12.575 1.130 12.825 1.270 ;
        RECT 11.595 0.880 12.825 1.130 ;
        RECT 11.595 0.365 11.910 0.880 ;
        RECT 12.575 0.350 12.825 0.880 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.440 3.415 ;
        RECT 0.110 2.520 0.360 3.245 ;
        RECT 0.560 2.520 0.890 2.980 ;
        RECT 1.090 2.650 1.340 3.245 ;
        RECT 2.005 2.680 2.335 3.245 ;
        RECT 0.685 2.480 0.890 2.520 ;
        RECT 3.030 2.510 3.360 2.755 ;
        RECT 1.510 2.480 3.360 2.510 ;
        RECT 0.685 2.340 3.360 2.480 ;
        RECT 3.560 2.570 3.810 2.755 ;
        RECT 4.400 2.740 4.730 3.245 ;
        RECT 4.915 2.570 5.180 2.755 ;
        RECT 5.830 2.745 6.165 3.245 ;
        RECT 3.560 2.400 5.180 2.570 ;
        RECT 0.685 2.310 1.680 2.340 ;
        RECT 0.685 0.830 0.855 2.310 ;
        RECT 3.030 2.230 3.360 2.340 ;
        RECT 1.025 1.130 1.285 2.140 ;
        RECT 1.455 1.810 1.805 2.140 ;
        RECT 2.455 1.890 2.845 2.170 ;
        RECT 3.030 2.060 3.795 2.230 ;
        RECT 1.455 1.140 1.625 1.810 ;
        RECT 2.455 1.720 3.455 1.890 ;
        RECT 2.445 1.140 2.675 1.550 ;
        RECT 1.455 0.970 2.675 1.140 ;
        RECT 0.165 0.660 0.855 0.830 ;
        RECT 0.165 0.370 0.495 0.660 ;
        RECT 1.065 0.085 1.235 0.830 ;
        RECT 1.455 0.350 1.875 0.970 ;
        RECT 2.845 0.800 3.015 1.720 ;
        RECT 3.190 1.560 3.455 1.720 ;
        RECT 3.625 1.390 3.795 2.060 ;
        RECT 2.045 0.085 2.375 0.800 ;
        RECT 2.545 0.500 3.015 0.800 ;
        RECT 3.185 1.220 3.795 1.390 ;
        RECT 3.185 0.670 3.435 1.220 ;
        RECT 3.965 1.050 4.135 2.400 ;
        RECT 4.745 2.295 5.180 2.400 ;
        RECT 5.395 2.405 6.955 2.575 ;
        RECT 7.125 2.475 8.410 2.805 ;
        RECT 3.605 0.880 4.135 1.050 ;
        RECT 4.305 1.050 4.570 2.105 ;
        RECT 4.745 1.500 4.915 2.295 ;
        RECT 5.395 2.290 5.725 2.405 ;
        RECT 5.085 1.670 5.635 2.120 ;
        RECT 6.155 1.940 6.615 2.235 ;
        RECT 4.745 1.220 5.985 1.500 ;
        RECT 6.155 1.050 6.325 1.940 ;
        RECT 6.785 1.590 6.955 2.405 ;
        RECT 6.495 1.260 6.955 1.590 ;
        RECT 4.305 0.880 6.990 1.050 ;
        RECT 3.605 0.670 3.935 0.880 ;
        RECT 5.735 0.720 6.990 0.880 ;
        RECT 7.160 0.845 7.330 2.475 ;
        RECT 7.740 1.345 8.070 2.305 ;
        RECT 8.240 1.705 8.410 2.475 ;
        RECT 8.580 2.445 8.910 3.245 ;
        RECT 9.080 2.445 9.480 2.905 ;
        RECT 9.650 2.445 9.900 3.245 ;
        RECT 8.765 1.920 9.140 2.275 ;
        RECT 9.310 2.045 9.480 2.445 ;
        RECT 9.310 1.875 9.945 2.045 ;
        RECT 8.240 1.535 9.605 1.705 ;
        RECT 9.345 1.375 9.605 1.535 ;
        RECT 7.545 1.015 8.275 1.345 ;
        RECT 8.445 1.205 8.775 1.365 ;
        RECT 9.775 1.205 9.945 1.875 ;
        RECT 10.115 1.630 10.365 2.905 ;
        RECT 10.535 2.025 10.865 3.245 ;
        RECT 11.535 2.140 12.240 3.245 ;
        RECT 12.910 1.950 13.240 3.245 ;
        RECT 10.115 1.460 12.240 1.630 ;
        RECT 8.445 1.035 9.945 1.205 ;
        RECT 10.560 1.300 12.240 1.460 ;
        RECT 4.305 0.540 5.565 0.710 ;
        RECT 7.160 0.595 7.935 0.845 ;
        RECT 4.305 0.500 4.475 0.540 ;
        RECT 2.545 0.330 4.475 0.500 ;
        RECT 5.395 0.425 5.565 0.540 ;
        RECT 8.105 0.425 8.275 1.015 ;
        RECT 4.895 0.085 5.225 0.370 ;
        RECT 5.395 0.255 8.275 0.425 ;
        RECT 8.625 0.085 8.955 0.845 ;
        RECT 9.500 0.385 9.830 1.035 ;
        RECT 10.115 0.085 10.390 1.130 ;
        RECT 10.560 0.350 10.890 1.300 ;
        RECT 11.120 0.085 11.410 1.130 ;
        RECT 12.080 0.085 12.405 0.710 ;
        RECT 13.005 0.085 13.335 1.100 ;
        RECT 0.000 -0.085 13.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 8.795 1.950 8.965 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
  END
END sky130_fd_sc_hs__dfrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.180 1.795 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.475 1.010 0.805 2.020 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.735 5.665 1.780 ;
        RECT 8.255 1.735 8.545 1.780 ;
        RECT 5.375 1.595 8.545 1.735 ;
        RECT 5.375 1.550 5.665 1.595 ;
        RECT 8.255 1.550 8.545 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.000 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 0.955 2.405 1.240 ;
        RECT 0.995 0.950 4.545 0.955 ;
        RECT 0.005 0.920 4.545 0.950 ;
        RECT 5.745 0.920 7.215 1.140 ;
        RECT 9.375 0.920 11.995 1.240 ;
        RECT 0.005 0.245 11.995 0.920 ;
        RECT 0.000 0.000 12.000 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 12.190 3.520 ;
        RECT 0.965 1.610 6.715 1.660 ;
        RECT 5.675 1.525 6.715 1.610 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.000 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 11.555 1.820 11.885 2.980 ;
        RECT 11.715 1.050 11.885 1.820 ;
        RECT 11.555 0.350 11.885 1.050 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 10.120 1.180 10.435 2.980 ;
        RECT 10.120 1.130 10.315 1.180 ;
        RECT 9.985 0.350 10.315 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.000 3.415 ;
        RECT 0.115 2.360 0.365 2.980 ;
        RECT 0.565 2.590 0.895 3.245 ;
        RECT 1.575 2.530 1.905 3.245 ;
        RECT 2.105 2.905 3.875 3.075 ;
        RECT 2.105 2.400 2.355 2.905 ;
        RECT 0.115 2.230 1.795 2.360 ;
        RECT 2.525 2.295 3.005 2.735 ;
        RECT 3.175 2.295 3.535 2.735 ;
        RECT 2.525 2.230 2.695 2.295 ;
        RECT 0.115 2.190 2.695 2.230 ;
        RECT 0.115 0.840 0.285 2.190 ;
        RECT 1.625 2.060 2.695 2.190 ;
        RECT 0.975 1.890 1.455 2.020 ;
        RECT 0.975 1.720 2.355 1.890 ;
        RECT 0.975 1.010 1.145 1.720 ;
        RECT 2.025 1.300 2.355 1.720 ;
        RECT 0.115 0.380 0.365 0.840 ;
        RECT 0.545 0.085 0.795 0.840 ;
        RECT 0.975 0.350 1.435 1.010 ;
        RECT 1.605 0.085 1.865 1.010 ;
        RECT 2.045 0.425 2.295 1.130 ;
        RECT 2.525 0.845 2.695 2.060 ;
        RECT 2.865 1.435 3.195 2.105 ;
        RECT 2.525 0.595 2.855 0.845 ;
        RECT 3.025 0.425 3.195 1.435 ;
        RECT 2.045 0.255 3.195 0.425 ;
        RECT 3.365 1.055 3.535 2.295 ;
        RECT 3.705 2.335 3.875 2.905 ;
        RECT 4.045 2.505 4.440 3.245 ;
        RECT 4.610 2.905 5.540 3.075 ;
        RECT 4.610 2.335 4.780 2.905 ;
        RECT 3.705 2.165 4.780 2.335 ;
        RECT 3.705 1.360 3.945 2.165 ;
        RECT 4.950 1.995 5.200 2.735 ;
        RECT 5.370 2.295 5.540 2.905 ;
        RECT 5.710 2.465 6.050 3.245 ;
        RECT 6.760 2.650 7.450 2.905 ;
        RECT 8.070 2.650 8.240 3.245 ;
        RECT 6.760 2.480 7.900 2.650 ;
        RECT 8.440 2.480 8.770 2.980 ;
        RECT 5.370 2.125 6.035 2.295 ;
        RECT 4.230 1.775 5.200 1.995 ;
        RECT 4.115 1.435 5.235 1.605 ;
        RECT 5.405 1.550 5.695 1.955 ;
        RECT 5.865 1.790 6.035 2.125 ;
        RECT 6.760 1.960 7.010 2.480 ;
        RECT 7.230 2.020 7.560 2.310 ;
        RECT 7.730 2.220 8.770 2.480 ;
        RECT 9.000 2.560 9.330 2.980 ;
        RECT 9.560 2.730 9.910 3.245 ;
        RECT 9.000 2.390 9.735 2.560 ;
        RECT 7.730 2.050 9.395 2.220 ;
        RECT 6.840 1.850 7.010 1.960 ;
        RECT 5.865 1.620 6.605 1.790 ;
        RECT 6.840 1.680 7.220 1.850 ;
        RECT 6.435 1.450 6.605 1.620 ;
        RECT 4.115 1.055 4.285 1.435 ;
        RECT 4.950 1.290 5.235 1.435 ;
        RECT 5.935 1.290 6.265 1.450 ;
        RECT 3.365 0.885 4.285 1.055 ;
        RECT 4.455 0.885 4.775 1.265 ;
        RECT 4.950 1.120 6.265 1.290 ;
        RECT 6.435 1.120 6.880 1.450 ;
        RECT 4.950 1.055 5.235 1.120 ;
        RECT 3.365 0.385 3.615 0.885 ;
        RECT 4.105 0.085 4.435 0.715 ;
        RECT 4.605 0.435 5.180 0.885 ;
        RECT 5.855 0.085 6.185 0.950 ;
        RECT 6.435 0.425 6.605 1.120 ;
        RECT 7.050 0.925 7.220 1.680 ;
        RECT 6.775 0.595 7.220 0.925 ;
        RECT 7.390 0.425 7.560 2.020 ;
        RECT 7.770 1.010 8.100 1.880 ;
        RECT 8.285 1.180 8.670 1.780 ;
        RECT 9.065 1.210 9.395 2.050 ;
        RECT 9.565 1.010 9.735 2.390 ;
        RECT 7.770 0.840 9.735 1.010 ;
        RECT 10.680 1.550 10.850 2.875 ;
        RECT 11.050 1.995 11.380 3.245 ;
        RECT 10.680 1.220 11.540 1.550 ;
        RECT 10.680 0.940 10.875 1.220 ;
        RECT 6.435 0.255 7.560 0.425 ;
        RECT 8.065 0.085 8.755 0.670 ;
        RECT 8.925 0.415 9.255 0.840 ;
        RECT 9.485 0.085 9.815 0.670 ;
        RECT 10.545 0.350 10.875 0.940 ;
        RECT 11.055 0.085 11.385 0.940 ;
        RECT 0.000 -0.085 12.000 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 5.435 1.580 5.605 1.750 ;
        RECT 8.315 1.580 8.485 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
  END
END sky130_fd_sc_hs__dfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfsbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.180 1.775 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.980 0.805 1.990 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.735 5.665 1.780 ;
        RECT 8.255 1.735 8.545 1.780 ;
        RECT 5.375 1.595 8.545 1.735 ;
        RECT 5.375 1.550 5.665 1.595 ;
        RECT 8.255 1.550 8.545 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.035 2.400 1.240 ;
        RECT 9.555 1.140 12.955 1.240 ;
        RECT 0.995 0.920 4.430 1.035 ;
        RECT 5.775 0.920 12.955 1.140 ;
        RECT 0.005 0.245 12.955 0.920 ;
        RECT 0.000 0.000 12.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.150 3.520 ;
        RECT 0.965 1.610 6.735 1.660 ;
        RECT 5.695 1.525 6.735 1.610 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.960 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 12.065 1.820 12.425 2.980 ;
        RECT 12.255 1.130 12.425 1.820 ;
        RECT 12.085 0.350 12.425 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 10.130 1.820 10.435 2.970 ;
        RECT 10.175 0.350 10.435 1.820 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.115 2.360 0.365 2.980 ;
        RECT 0.565 2.530 0.895 3.245 ;
        RECT 1.575 2.530 1.905 3.245 ;
        RECT 2.105 2.905 3.845 3.075 ;
        RECT 2.105 2.400 2.275 2.905 ;
        RECT 0.115 2.230 1.795 2.360 ;
        RECT 2.445 2.295 2.865 2.735 ;
        RECT 3.065 2.295 3.455 2.735 ;
        RECT 2.445 2.230 2.615 2.295 ;
        RECT 0.115 2.190 2.615 2.230 ;
        RECT 0.115 0.810 0.285 2.190 ;
        RECT 1.625 2.060 2.615 2.190 ;
        RECT 0.975 1.890 1.455 2.020 ;
        RECT 0.975 1.720 2.275 1.890 ;
        RECT 0.975 1.010 1.145 1.720 ;
        RECT 1.945 1.300 2.275 1.720 ;
        RECT 0.115 0.350 0.365 0.810 ;
        RECT 0.545 0.085 0.795 0.810 ;
        RECT 0.975 0.350 1.435 1.010 ;
        RECT 1.605 0.085 1.865 1.010 ;
        RECT 2.045 0.425 2.215 1.130 ;
        RECT 2.445 0.925 2.615 2.060 ;
        RECT 2.785 1.435 3.115 2.105 ;
        RECT 2.445 0.595 2.770 0.925 ;
        RECT 2.940 0.425 3.110 1.435 ;
        RECT 3.285 1.265 3.455 2.295 ;
        RECT 3.625 2.565 3.845 2.905 ;
        RECT 4.020 2.735 4.350 3.245 ;
        RECT 4.520 2.905 5.530 3.075 ;
        RECT 4.520 2.565 4.690 2.905 ;
        RECT 3.625 2.395 4.690 2.565 ;
        RECT 3.625 1.435 3.845 2.395 ;
        RECT 4.860 2.295 5.190 2.735 ;
        RECT 5.360 2.360 5.530 2.905 ;
        RECT 5.700 2.530 6.070 3.245 ;
        RECT 6.780 2.650 7.470 2.980 ;
        RECT 8.090 2.650 8.260 3.245 ;
        RECT 6.780 2.480 7.920 2.650 ;
        RECT 8.460 2.480 8.790 2.915 ;
        RECT 9.630 2.630 9.960 3.245 ;
        RECT 4.860 2.225 5.030 2.295 ;
        RECT 4.140 2.055 5.030 2.225 ;
        RECT 5.360 2.190 6.500 2.360 ;
        RECT 4.140 1.855 4.470 2.055 ;
        RECT 4.750 1.685 5.015 1.885 ;
        RECT 4.015 1.515 5.015 1.685 ;
        RECT 5.225 1.580 5.635 2.020 ;
        RECT 4.015 1.265 4.185 1.515 ;
        RECT 4.750 1.410 5.015 1.515 ;
        RECT 6.330 1.450 6.500 2.190 ;
        RECT 6.780 1.850 7.030 2.480 ;
        RECT 7.250 2.020 7.580 2.310 ;
        RECT 7.750 2.120 8.790 2.480 ;
        RECT 9.015 2.460 9.345 2.620 ;
        RECT 9.015 2.290 9.910 2.460 ;
        RECT 6.780 1.680 7.215 1.850 ;
        RECT 3.285 1.095 4.185 1.265 ;
        RECT 3.285 0.925 3.530 1.095 ;
        RECT 4.355 1.015 4.580 1.345 ;
        RECT 4.750 1.240 5.915 1.410 ;
        RECT 5.585 1.120 5.915 1.240 ;
        RECT 6.330 1.120 6.875 1.450 ;
        RECT 3.280 0.465 3.530 0.925 ;
        RECT 2.045 0.255 3.110 0.425 ;
        RECT 3.990 0.085 4.240 0.845 ;
        RECT 4.410 0.350 4.880 1.015 ;
        RECT 5.340 0.085 6.160 0.680 ;
        RECT 6.330 0.450 6.500 1.120 ;
        RECT 7.045 0.950 7.215 1.680 ;
        RECT 6.670 0.620 7.215 0.950 ;
        RECT 7.385 0.450 7.555 2.020 ;
        RECT 7.750 1.950 9.570 2.120 ;
        RECT 7.725 1.010 8.055 1.780 ;
        RECT 8.285 1.180 8.640 1.780 ;
        RECT 8.900 1.350 9.570 1.950 ;
        RECT 9.740 1.180 9.910 2.290 ;
        RECT 10.605 1.820 10.860 3.245 ;
        RECT 9.105 1.010 9.910 1.180 ;
        RECT 11.085 1.630 11.415 2.860 ;
        RECT 11.615 1.820 11.865 3.245 ;
        RECT 12.595 1.820 12.845 3.245 ;
        RECT 11.085 1.300 12.085 1.630 ;
        RECT 7.725 0.840 9.435 1.010 ;
        RECT 6.330 0.280 7.555 0.450 ;
        RECT 8.100 0.085 8.845 0.670 ;
        RECT 9.105 0.635 9.435 0.840 ;
        RECT 9.665 0.085 9.995 0.840 ;
        RECT 10.605 0.085 10.855 1.130 ;
        RECT 11.085 0.350 11.415 1.300 ;
        RECT 11.585 0.085 11.915 1.030 ;
        RECT 12.595 0.085 12.845 1.130 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 5.435 1.580 5.605 1.750 ;
        RECT 8.315 1.580 8.485 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
  END
END sky130_fd_sc_hs__dfsbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.180 1.795 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.980 0.805 1.990 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 8.255 2.105 8.545 2.150 ;
        RECT 5.375 1.965 8.545 2.105 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 8.255 1.920 8.545 1.965 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.035 2.385 1.240 ;
        RECT 0.995 0.920 2.925 1.035 ;
        RECT 4.575 0.920 7.015 1.140 ;
        RECT 9.890 1.050 10.940 1.240 ;
        RECT 9.380 0.920 10.940 1.050 ;
        RECT 0.005 0.245 10.940 0.920 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
        RECT 0.940 1.570 6.430 1.660 ;
        RECT 5.390 1.525 6.430 1.570 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.050 10.935 2.980 ;
        RECT 10.500 0.350 10.935 1.050 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.105 2.400 0.355 2.980 ;
        RECT 0.555 2.570 0.885 3.245 ;
        RECT 1.540 2.570 1.870 3.245 ;
        RECT 2.070 2.905 3.755 3.075 ;
        RECT 2.070 2.400 2.320 2.905 ;
        RECT 0.105 2.230 1.760 2.400 ;
        RECT 2.490 2.295 2.910 2.735 ;
        RECT 3.080 2.295 3.415 2.735 ;
        RECT 2.490 2.230 2.660 2.295 ;
        RECT 0.105 0.810 0.275 2.230 ;
        RECT 1.590 2.060 2.660 2.230 ;
        RECT 0.975 1.890 1.420 2.060 ;
        RECT 0.975 1.720 2.315 1.890 ;
        RECT 0.975 1.010 1.145 1.720 ;
        RECT 1.985 1.260 2.315 1.720 ;
        RECT 0.105 0.350 0.365 0.810 ;
        RECT 0.545 0.085 0.795 0.810 ;
        RECT 0.975 0.350 1.435 1.010 ;
        RECT 1.615 0.085 1.785 1.010 ;
        RECT 1.965 0.425 2.295 1.090 ;
        RECT 2.485 0.925 2.660 2.060 ;
        RECT 2.830 1.435 3.075 2.105 ;
        RECT 2.485 0.595 2.735 0.925 ;
        RECT 2.905 0.425 3.075 1.435 ;
        RECT 1.965 0.255 3.075 0.425 ;
        RECT 3.245 1.020 3.415 2.295 ;
        RECT 3.585 2.255 3.755 2.905 ;
        RECT 3.950 2.425 4.230 3.245 ;
        RECT 4.400 2.905 5.365 3.075 ;
        RECT 4.400 2.255 4.570 2.905 ;
        RECT 3.585 2.085 4.570 2.255 ;
        RECT 4.740 2.320 5.025 2.735 ;
        RECT 5.195 2.490 5.365 2.905 ;
        RECT 5.535 2.660 5.785 3.245 ;
        RECT 6.475 2.625 7.600 2.980 ;
        RECT 7.770 2.650 7.940 3.245 ;
        RECT 5.195 2.320 5.975 2.490 ;
        RECT 3.585 1.435 3.755 2.085 ;
        RECT 4.740 1.915 4.910 2.320 ;
        RECT 4.055 1.745 4.910 1.915 ;
        RECT 5.080 1.820 5.635 2.150 ;
        RECT 5.805 1.885 5.975 2.320 ;
        RECT 6.475 2.050 6.810 2.625 ;
        RECT 7.430 2.480 7.600 2.625 ;
        RECT 8.140 2.480 8.470 2.930 ;
        RECT 8.665 2.650 8.915 3.245 ;
        RECT 9.115 2.650 9.445 2.980 ;
        RECT 4.055 1.685 4.385 1.745 ;
        RECT 5.805 1.715 6.405 1.885 ;
        RECT 4.805 1.515 6.065 1.545 ;
        RECT 3.925 1.345 6.065 1.515 ;
        RECT 3.925 1.020 4.095 1.345 ;
        RECT 4.805 1.215 6.065 1.345 ;
        RECT 6.235 1.450 6.405 1.715 ;
        RECT 6.575 1.800 6.810 2.050 ;
        RECT 6.980 2.140 7.260 2.355 ;
        RECT 7.430 2.310 9.105 2.480 ;
        RECT 6.980 1.970 7.325 2.140 ;
        RECT 6.575 1.630 6.985 1.800 ;
        RECT 3.245 0.850 4.095 1.020 ;
        RECT 4.265 1.030 4.625 1.175 ;
        RECT 6.235 1.120 6.645 1.450 ;
        RECT 4.265 0.860 5.010 1.030 ;
        RECT 3.245 0.415 3.575 0.850 ;
        RECT 4.065 0.085 4.455 0.680 ;
        RECT 4.625 0.570 5.010 0.860 ;
        RECT 5.620 0.085 5.950 1.030 ;
        RECT 6.235 0.425 6.405 1.120 ;
        RECT 6.815 0.925 6.985 1.630 ;
        RECT 6.575 0.595 6.985 0.925 ;
        RECT 7.155 0.425 7.325 1.970 ;
        RECT 7.495 0.960 7.730 1.555 ;
        RECT 8.185 1.130 8.515 2.140 ;
        RECT 8.775 1.370 9.105 2.310 ;
        RECT 9.275 1.200 9.445 2.650 ;
        RECT 9.090 1.030 9.445 1.200 ;
        RECT 9.635 1.550 9.965 2.875 ;
        RECT 10.155 1.820 10.485 3.245 ;
        RECT 9.635 1.220 10.515 1.550 ;
        RECT 9.090 0.960 9.260 1.030 ;
        RECT 7.495 0.790 9.260 0.960 ;
        RECT 9.635 0.860 9.820 1.220 ;
        RECT 6.235 0.255 7.325 0.425 ;
        RECT 7.870 0.085 8.760 0.600 ;
        RECT 8.930 0.350 9.260 0.790 ;
        RECT 9.490 0.350 9.820 0.860 ;
        RECT 10.000 0.085 10.330 1.030 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 8.315 1.950 8.485 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__dfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfstp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.180 1.775 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.980 0.805 1.990 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 5.855 2.105 6.145 2.150 ;
        RECT 8.255 2.105 8.545 2.150 ;
        RECT 5.855 1.965 8.545 2.105 ;
        RECT 5.855 1.920 6.145 1.965 ;
        RECT 8.255 1.920 8.545 1.965 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.000 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.035 2.405 1.240 ;
        RECT 9.980 1.140 11.995 1.240 ;
        RECT 0.995 0.920 2.965 1.035 ;
        RECT 4.720 0.920 11.995 1.140 ;
        RECT 0.005 0.245 11.995 0.920 ;
        RECT 0.000 0.000 12.000 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 12.190 3.520 ;
        RECT 0.965 1.610 6.775 1.660 ;
        RECT 5.735 1.525 6.775 1.610 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.000 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 11.155 2.150 11.465 2.980 ;
        RECT 10.685 1.820 11.465 2.150 ;
        RECT 11.295 1.130 11.465 1.820 ;
        RECT 11.100 0.350 11.465 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.000 3.415 ;
        RECT 0.115 2.360 0.365 2.980 ;
        RECT 0.565 2.530 0.895 3.245 ;
        RECT 1.575 2.530 1.905 3.245 ;
        RECT 2.105 2.890 3.795 3.060 ;
        RECT 2.105 2.400 2.275 2.890 ;
        RECT 0.115 2.230 1.795 2.360 ;
        RECT 2.445 2.260 2.945 2.720 ;
        RECT 3.115 2.260 3.455 2.720 ;
        RECT 2.445 2.230 2.615 2.260 ;
        RECT 0.115 2.190 2.615 2.230 ;
        RECT 0.115 0.765 0.285 2.190 ;
        RECT 1.625 2.060 2.615 2.190 ;
        RECT 0.975 1.890 1.455 2.020 ;
        RECT 0.975 1.720 2.275 1.890 ;
        RECT 0.975 1.010 1.145 1.720 ;
        RECT 1.945 1.300 2.275 1.720 ;
        RECT 0.115 0.395 0.365 0.765 ;
        RECT 0.545 0.085 0.795 0.765 ;
        RECT 0.975 0.350 1.435 1.010 ;
        RECT 1.615 0.085 1.865 1.010 ;
        RECT 2.045 0.425 2.215 1.130 ;
        RECT 2.445 0.925 2.615 2.060 ;
        RECT 2.785 1.380 3.115 2.050 ;
        RECT 2.445 0.595 2.775 0.925 ;
        RECT 2.945 0.425 3.115 1.380 ;
        RECT 2.045 0.255 3.115 0.425 ;
        RECT 3.285 1.210 3.455 2.260 ;
        RECT 3.625 2.410 3.795 2.890 ;
        RECT 4.070 2.910 4.240 3.245 ;
        RECT 4.070 2.580 4.575 2.910 ;
        RECT 4.745 2.890 5.690 3.060 ;
        RECT 4.745 2.410 4.915 2.890 ;
        RECT 3.625 2.240 4.915 2.410 ;
        RECT 5.085 2.320 5.350 2.720 ;
        RECT 5.520 2.490 5.690 2.890 ;
        RECT 5.860 2.660 6.110 3.245 ;
        RECT 6.820 2.730 7.470 2.980 ;
        RECT 6.820 2.550 7.930 2.730 ;
        RECT 8.100 2.720 8.430 3.245 ;
        RECT 8.630 2.550 8.880 2.980 ;
        RECT 9.110 2.660 9.440 3.245 ;
        RECT 5.520 2.320 6.585 2.490 ;
        RECT 3.625 1.380 3.915 2.240 ;
        RECT 5.085 2.070 5.255 2.320 ;
        RECT 4.230 1.740 5.255 2.070 ;
        RECT 5.425 1.790 6.115 2.150 ;
        RECT 4.085 1.400 6.245 1.570 ;
        RECT 4.085 1.210 4.255 1.400 ;
        RECT 3.285 1.040 4.255 1.210 ;
        RECT 4.425 1.050 4.770 1.230 ;
        RECT 4.950 1.220 6.245 1.400 ;
        RECT 5.915 1.215 6.245 1.220 ;
        RECT 6.415 1.450 6.585 2.320 ;
        RECT 6.820 1.790 7.070 2.550 ;
        RECT 7.760 2.490 8.880 2.550 ;
        RECT 7.290 2.150 7.590 2.380 ;
        RECT 7.760 2.320 9.470 2.490 ;
        RECT 7.290 1.980 7.660 2.150 ;
        RECT 6.820 1.620 7.320 1.790 ;
        RECT 6.415 1.120 6.960 1.450 ;
        RECT 3.285 0.400 3.615 1.040 ;
        RECT 4.425 0.880 5.160 1.050 ;
        RECT 4.270 0.085 4.600 0.710 ;
        RECT 4.770 0.570 5.160 0.880 ;
        RECT 5.650 0.085 6.245 1.030 ;
        RECT 6.415 0.450 6.585 1.120 ;
        RECT 7.150 0.950 7.320 1.620 ;
        RECT 6.825 0.620 7.320 0.950 ;
        RECT 7.490 0.450 7.660 1.980 ;
        RECT 7.830 1.240 8.145 2.130 ;
        RECT 8.315 1.480 8.730 2.150 ;
        RECT 9.140 1.615 9.470 2.320 ;
        RECT 9.640 1.240 9.890 2.980 ;
        RECT 7.830 1.070 9.890 1.240 ;
        RECT 6.415 0.280 7.660 0.450 ;
        RECT 8.525 0.085 9.360 0.900 ;
        RECT 9.530 0.635 9.890 1.070 ;
        RECT 10.090 1.630 10.450 2.860 ;
        RECT 10.655 2.320 10.985 3.245 ;
        RECT 11.635 1.820 11.885 3.245 ;
        RECT 10.090 1.300 11.125 1.630 ;
        RECT 10.090 0.450 10.420 1.300 ;
        RECT 10.600 0.085 10.930 1.130 ;
        RECT 11.635 0.085 11.885 1.130 ;
        RECT 0.000 -0.085 12.000 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 5.915 1.950 6.085 2.120 ;
        RECT 8.315 1.950 8.485 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
  END
END sky130_fd_sc_hs__dfstp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfstp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.180 1.775 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.980 0.805 1.990 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.735 5.665 1.780 ;
        RECT 8.255 1.735 8.545 1.780 ;
        RECT 5.375 1.595 8.545 1.735 ;
        RECT 5.375 1.550 5.665 1.595 ;
        RECT 8.255 1.550 8.545 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.035 2.405 1.240 ;
        RECT 0.995 0.920 2.965 1.035 ;
        RECT 4.540 0.990 7.085 1.140 ;
        RECT 9.570 0.990 12.955 1.240 ;
        RECT 4.540 0.920 12.955 0.990 ;
        RECT 0.005 0.245 12.955 0.920 ;
        RECT 0.000 0.000 12.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.150 3.520 ;
        RECT 5.505 1.555 6.545 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.960 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.119700 ;
    PORT
      LAYER li1 ;
        RECT 11.175 2.080 11.455 2.980 ;
        RECT 12.125 2.150 12.355 2.980 ;
        RECT 12.125 2.080 12.835 2.150 ;
        RECT 11.175 1.820 12.835 2.080 ;
        RECT 12.605 1.150 12.835 1.820 ;
        RECT 10.680 0.980 12.835 1.150 ;
        RECT 10.680 0.350 11.010 0.980 ;
        RECT 12.015 0.350 12.345 0.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.115 2.410 0.365 2.960 ;
        RECT 0.565 2.580 0.895 3.245 ;
        RECT 1.575 2.580 1.905 3.245 ;
        RECT 2.105 2.905 3.795 3.075 ;
        RECT 2.105 2.410 2.275 2.905 ;
        RECT 0.115 2.240 1.795 2.410 ;
        RECT 2.445 2.295 2.945 2.735 ;
        RECT 3.115 2.295 3.455 2.735 ;
        RECT 2.445 2.240 2.615 2.295 ;
        RECT 0.115 0.810 0.285 2.240 ;
        RECT 1.625 2.070 2.615 2.240 ;
        RECT 0.975 1.890 1.455 2.070 ;
        RECT 0.975 1.720 2.275 1.890 ;
        RECT 0.975 1.010 1.145 1.720 ;
        RECT 1.945 1.350 2.275 1.720 ;
        RECT 0.115 0.350 0.365 0.810 ;
        RECT 0.545 0.085 0.795 0.810 ;
        RECT 0.975 0.340 1.435 1.010 ;
        RECT 1.615 0.085 1.865 1.010 ;
        RECT 2.045 0.425 2.215 1.130 ;
        RECT 2.445 0.925 2.615 2.070 ;
        RECT 2.785 1.455 3.115 2.125 ;
        RECT 2.445 0.595 2.775 0.925 ;
        RECT 2.945 0.425 3.115 1.455 ;
        RECT 2.045 0.255 3.115 0.425 ;
        RECT 3.285 1.300 3.455 2.295 ;
        RECT 3.625 2.335 3.795 2.905 ;
        RECT 3.985 2.755 4.155 3.245 ;
        RECT 4.515 2.905 5.510 3.075 ;
        RECT 3.985 2.505 4.345 2.755 ;
        RECT 4.515 2.335 4.685 2.905 ;
        RECT 3.625 2.165 4.685 2.335 ;
        RECT 4.855 2.295 5.170 2.735 ;
        RECT 3.625 1.470 3.795 2.165 ;
        RECT 4.855 1.995 5.025 2.295 ;
        RECT 5.340 2.265 5.510 2.905 ;
        RECT 5.680 2.435 5.940 3.245 ;
        RECT 6.590 2.650 7.265 2.980 ;
        RECT 7.885 2.650 8.055 3.245 ;
        RECT 6.670 2.480 7.715 2.650 ;
        RECT 8.255 2.480 8.585 2.980 ;
        RECT 8.780 2.650 9.030 3.245 ;
        RECT 9.230 2.650 9.560 2.980 ;
        RECT 5.340 2.095 6.475 2.265 ;
        RECT 4.115 1.740 5.025 1.995 ;
        RECT 3.965 1.400 5.025 1.570 ;
        RECT 5.195 1.550 5.635 1.925 ;
        RECT 3.965 1.300 4.135 1.400 ;
        RECT 3.285 1.130 4.135 1.300 ;
        RECT 4.770 1.370 5.025 1.400 ;
        RECT 5.805 1.370 6.135 1.490 ;
        RECT 3.285 0.350 3.535 1.130 ;
        RECT 4.305 0.950 4.590 1.230 ;
        RECT 4.770 1.200 6.135 1.370 ;
        RECT 6.305 1.450 6.475 2.095 ;
        RECT 6.670 1.790 6.840 2.480 ;
        RECT 7.545 2.310 9.110 2.480 ;
        RECT 7.045 2.020 7.375 2.310 ;
        RECT 6.670 1.620 7.035 1.790 ;
        RECT 4.770 1.120 5.025 1.200 ;
        RECT 6.305 1.120 6.695 1.450 ;
        RECT 4.305 0.780 5.050 0.950 ;
        RECT 4.590 0.620 5.050 0.780 ;
        RECT 4.025 0.085 4.420 0.600 ;
        RECT 5.670 0.085 6.000 1.030 ;
        RECT 6.305 0.425 6.475 1.120 ;
        RECT 6.865 0.925 7.035 1.620 ;
        RECT 6.645 0.595 7.035 0.925 ;
        RECT 7.205 0.425 7.375 2.020 ;
        RECT 7.545 1.010 7.875 1.655 ;
        RECT 8.185 1.180 8.515 1.850 ;
        RECT 8.780 1.370 9.110 2.310 ;
        RECT 9.280 1.010 9.450 2.650 ;
        RECT 9.755 1.820 10.005 3.245 ;
        RECT 10.205 1.650 10.535 2.700 ;
        RECT 10.725 1.820 11.005 3.245 ;
        RECT 11.625 2.250 11.955 3.245 ;
        RECT 12.525 2.320 12.855 3.245 ;
        RECT 10.205 1.490 11.995 1.650 ;
        RECT 7.545 0.840 9.450 1.010 ;
        RECT 6.305 0.255 7.375 0.425 ;
        RECT 7.935 0.085 8.950 0.670 ;
        RECT 9.120 0.420 9.450 0.840 ;
        RECT 9.680 1.320 11.995 1.490 ;
        RECT 9.680 0.350 10.010 1.320 ;
        RECT 10.180 0.085 10.510 1.130 ;
        RECT 11.180 0.085 11.845 0.800 ;
        RECT 12.515 0.085 12.845 0.810 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 5.435 1.580 5.605 1.750 ;
        RECT 8.315 1.580 8.485 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
  END
END sky130_fd_sc_hs__dfstp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.500 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.700 2.025 2.080 2.355 ;
        RECT 1.910 1.780 2.080 2.025 ;
        RECT 1.910 1.125 2.270 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.155 1.240 1.705 1.430 ;
        RECT 0.005 1.145 1.705 1.240 ;
        RECT 4.460 1.240 6.520 1.280 ;
        RECT 0.005 1.060 3.470 1.145 ;
        RECT 4.460 1.060 9.580 1.240 ;
        RECT 0.005 0.245 9.580 1.060 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 7.665 2.030 8.070 2.980 ;
        RECT 7.900 1.130 8.070 2.030 ;
        RECT 7.640 0.350 8.070 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.535700 ;
    PORT
      LAYER li1 ;
        RECT 9.160 1.820 9.515 2.980 ;
        RECT 9.345 1.130 9.515 1.820 ;
        RECT 9.140 0.350 9.515 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.110 1.890 0.360 2.980 ;
        RECT 0.560 2.060 0.810 3.245 ;
        RECT 1.010 2.715 1.340 2.980 ;
        RECT 1.555 2.885 1.885 3.245 ;
        RECT 3.740 2.925 4.130 3.245 ;
        RECT 4.300 2.905 5.990 3.075 ;
        RECT 2.055 2.755 3.290 2.885 ;
        RECT 4.300 2.800 5.150 2.905 ;
        RECT 4.300 2.755 4.470 2.800 ;
        RECT 2.055 2.715 4.470 2.755 ;
        RECT 1.010 2.545 2.225 2.715 ;
        RECT 3.120 2.585 4.470 2.715 ;
        RECT 0.110 1.720 0.840 1.890 ;
        RECT 1.010 1.815 1.435 2.545 ;
        RECT 2.780 2.415 2.950 2.545 ;
        RECT 2.250 2.045 2.610 2.375 ;
        RECT 0.670 1.550 0.840 1.720 ;
        RECT 0.115 0.900 0.445 1.010 ;
        RECT 0.670 0.900 1.090 1.550 ;
        RECT 1.265 1.485 1.740 1.815 ;
        RECT 1.265 1.070 1.595 1.485 ;
        RECT 2.440 1.240 2.610 2.045 ;
        RECT 2.780 2.245 4.280 2.415 ;
        RECT 2.780 1.580 2.950 2.245 ;
        RECT 3.120 1.750 3.655 2.075 ;
        RECT 2.780 1.410 3.315 1.580 ;
        RECT 2.440 1.070 2.885 1.240 ;
        RECT 0.115 0.730 2.545 0.900 ;
        RECT 0.115 0.350 0.445 0.730 ;
        RECT 0.625 0.085 1.005 0.560 ;
        RECT 1.855 0.085 2.205 0.560 ;
        RECT 2.375 0.425 2.545 0.730 ;
        RECT 2.715 0.595 2.885 1.070 ;
        RECT 3.065 0.595 3.315 1.410 ;
        RECT 3.485 0.750 3.655 1.750 ;
        RECT 4.020 1.630 4.280 2.245 ;
        RECT 4.640 2.025 4.810 2.615 ;
        RECT 4.450 1.855 4.810 2.025 ;
        RECT 4.450 1.370 4.620 1.855 ;
        RECT 4.980 1.685 5.150 2.800 ;
        RECT 3.825 1.185 4.620 1.370 ;
        RECT 4.790 1.355 5.150 1.685 ;
        RECT 5.320 2.115 5.570 2.735 ;
        RECT 5.320 1.380 5.490 2.115 ;
        RECT 5.820 1.945 5.990 2.905 ;
        RECT 6.165 2.390 6.495 3.245 ;
        RECT 6.710 2.220 7.040 2.860 ;
        RECT 5.660 1.615 5.990 1.945 ;
        RECT 6.230 1.860 7.040 2.220 ;
        RECT 7.240 2.030 7.490 3.245 ;
        RECT 6.230 1.690 7.730 1.860 ;
        RECT 6.230 1.550 6.560 1.690 ;
        RECT 6.800 1.380 7.130 1.520 ;
        RECT 5.320 1.210 7.130 1.380 ;
        RECT 3.825 1.015 4.900 1.185 ;
        RECT 5.320 1.120 5.590 1.210 ;
        RECT 6.800 1.190 7.130 1.210 ;
        RECT 7.300 1.350 7.730 1.690 ;
        RECT 8.280 1.630 8.455 2.700 ;
        RECT 8.655 1.820 8.985 3.245 ;
        RECT 4.570 0.920 4.900 1.015 ;
        RECT 5.125 0.790 5.590 1.120 ;
        RECT 3.485 0.620 4.650 0.750 ;
        RECT 3.485 0.580 5.715 0.620 ;
        RECT 3.485 0.425 3.655 0.580 ;
        RECT 2.375 0.255 3.655 0.425 ;
        RECT 3.980 0.085 4.310 0.410 ;
        RECT 4.480 0.290 5.715 0.580 ;
        RECT 6.080 0.085 6.410 1.040 ;
        RECT 7.300 1.020 7.470 1.350 ;
        RECT 6.640 0.850 7.470 1.020 ;
        RECT 8.280 1.300 9.175 1.630 ;
        RECT 6.640 0.440 6.970 0.850 ;
        RECT 7.140 0.085 7.470 0.680 ;
        RECT 8.280 0.625 8.530 1.300 ;
        RECT 8.710 0.085 8.960 1.130 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
  END
END sky130_fd_sc_hs__dfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.585 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.825 2.025 2.155 2.355 ;
        RECT 1.985 1.780 2.155 2.025 ;
        RECT 1.985 1.125 2.375 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.160 1.240 1.710 1.430 ;
        RECT 0.005 1.145 1.710 1.240 ;
        RECT 4.445 1.190 4.995 1.560 ;
        RECT 7.105 1.240 9.060 1.260 ;
        RECT 7.105 1.190 11.035 1.240 ;
        RECT 0.005 1.060 3.490 1.145 ;
        RECT 4.445 1.060 11.035 1.190 ;
        RECT 0.005 0.245 11.035 1.060 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.940 11.230 3.520 ;
        RECT -0.190 1.660 3.700 1.940 ;
        RECT 5.205 1.660 11.230 1.940 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 8.145 1.550 8.515 2.070 ;
        RECT 8.145 0.370 8.450 1.550 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 10.140 1.820 10.505 2.980 ;
        RECT 10.335 1.130 10.505 1.820 ;
        RECT 10.165 0.350 10.505 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.115 1.890 0.445 2.980 ;
        RECT 0.645 2.060 0.895 3.245 ;
        RECT 1.095 2.795 1.345 2.980 ;
        RECT 1.575 2.965 2.035 3.245 ;
        RECT 4.000 2.965 4.330 3.245 ;
        RECT 5.035 2.795 6.205 2.965 ;
        RECT 1.095 2.625 5.205 2.795 ;
        RECT 0.115 1.720 0.925 1.890 ;
        RECT 1.095 1.815 1.440 2.625 ;
        RECT 2.325 2.205 2.715 2.455 ;
        RECT 0.755 1.550 0.925 1.720 ;
        RECT 0.755 1.010 1.100 1.550 ;
        RECT 1.270 1.485 1.815 1.815 ;
        RECT 1.270 1.070 1.600 1.485 ;
        RECT 2.545 1.240 2.715 2.205 ;
        RECT 2.885 2.285 4.325 2.455 ;
        RECT 2.885 1.580 3.055 2.285 ;
        RECT 3.225 1.750 3.640 2.065 ;
        RECT 2.885 1.410 3.300 1.580 ;
        RECT 2.545 1.070 2.870 1.240 ;
        RECT 0.115 0.900 1.100 1.010 ;
        RECT 0.115 0.730 2.530 0.900 ;
        RECT 0.115 0.350 0.445 0.730 ;
        RECT 0.625 0.085 1.010 0.560 ;
        RECT 1.860 0.085 2.190 0.560 ;
        RECT 2.360 0.425 2.530 0.730 ;
        RECT 2.700 0.595 2.870 1.070 ;
        RECT 3.050 0.595 3.300 1.410 ;
        RECT 3.470 0.950 3.640 1.750 ;
        RECT 4.155 1.960 4.325 2.285 ;
        RECT 4.535 2.180 4.865 2.455 ;
        RECT 4.155 1.630 4.475 1.960 ;
        RECT 4.645 1.450 4.815 2.180 ;
        RECT 5.035 1.450 5.205 2.625 ;
        RECT 5.375 1.790 5.705 2.625 ;
        RECT 5.875 1.960 6.205 2.795 ;
        RECT 6.600 2.375 6.930 3.245 ;
        RECT 7.160 2.410 7.490 2.980 ;
        RECT 7.695 2.580 8.025 3.245 ;
        RECT 8.595 2.580 8.925 3.245 ;
        RECT 7.160 2.240 9.015 2.410 ;
        RECT 7.160 2.130 7.925 2.240 ;
        RECT 6.375 1.790 7.585 1.960 ;
        RECT 5.375 1.670 7.585 1.790 ;
        RECT 5.375 1.620 6.545 1.670 ;
        RECT 3.810 1.120 4.815 1.450 ;
        RECT 4.985 1.120 5.275 1.450 ;
        RECT 5.445 1.170 5.845 1.450 ;
        RECT 3.470 0.780 4.815 0.950 ;
        RECT 3.470 0.425 3.640 0.780 ;
        RECT 2.360 0.255 3.640 0.425 ;
        RECT 4.030 0.085 4.370 0.610 ;
        RECT 4.645 0.530 4.815 0.780 ;
        RECT 5.445 0.530 5.615 1.170 ;
        RECT 6.015 0.950 6.185 1.620 ;
        RECT 7.755 1.500 7.925 2.130 ;
        RECT 6.715 1.330 7.925 1.500 ;
        RECT 6.715 1.170 7.465 1.330 ;
        RECT 8.685 1.320 9.015 2.240 ;
        RECT 9.235 1.630 9.485 2.860 ;
        RECT 9.690 1.820 9.940 3.245 ;
        RECT 10.675 1.820 10.925 3.245 ;
        RECT 5.785 0.700 6.185 0.950 ;
        RECT 4.645 0.255 6.240 0.530 ;
        RECT 6.655 0.085 6.985 1.000 ;
        RECT 7.215 0.370 7.465 1.170 ;
        RECT 9.235 1.300 10.165 1.630 ;
        RECT 7.645 0.085 7.975 1.150 ;
        RECT 8.620 0.085 8.950 1.150 ;
        RECT 9.235 0.450 9.510 1.300 ;
        RECT 9.735 0.085 9.985 1.130 ;
        RECT 10.675 0.085 10.925 1.130 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__dfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.505 1.780 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.870 2.025 2.250 2.355 ;
        RECT 1.970 1.125 2.250 2.025 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.465 1.240 3.085 1.430 ;
        RECT 0.005 1.175 3.085 1.240 ;
        RECT 0.005 1.055 3.560 1.175 ;
        RECT 7.210 1.170 8.155 1.240 ;
        RECT 4.640 1.055 8.155 1.170 ;
        RECT 0.005 0.245 8.155 1.055 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 7.715 2.030 8.075 2.980 ;
        RECT 7.905 1.130 8.075 2.030 ;
        RECT 7.715 0.350 8.075 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.645 2.290 0.815 3.245 ;
        RECT 1.015 2.795 1.345 2.980 ;
        RECT 1.575 2.965 1.910 3.245 ;
        RECT 3.800 2.965 4.130 3.245 ;
        RECT 2.080 2.795 3.460 2.965 ;
        RECT 4.780 2.905 5.840 3.075 ;
        RECT 4.780 2.795 4.950 2.905 ;
        RECT 1.015 2.625 2.250 2.795 ;
        RECT 3.290 2.625 4.950 2.795 ;
        RECT 0.115 1.950 0.845 2.120 ;
        RECT 0.675 1.550 0.845 1.950 ;
        RECT 1.015 1.820 1.475 2.625 ;
        RECT 1.305 1.680 1.475 1.820 ;
        RECT 0.675 1.130 1.135 1.550 ;
        RECT 0.115 0.960 1.135 1.130 ;
        RECT 0.115 0.350 0.365 0.960 ;
        RECT 0.545 0.085 0.795 0.790 ;
        RECT 0.965 0.425 1.135 0.960 ;
        RECT 1.305 1.350 1.760 1.680 ;
        RECT 1.305 0.595 1.475 1.350 ;
        RECT 2.420 1.240 2.590 2.625 ;
        RECT 2.760 2.455 3.120 2.625 ;
        RECT 2.760 2.285 4.140 2.455 ;
        RECT 2.760 1.580 2.930 2.285 ;
        RECT 3.100 1.750 3.760 2.080 ;
        RECT 2.760 1.410 3.420 1.580 ;
        RECT 2.420 1.070 2.975 1.240 ;
        RECT 1.645 0.730 2.655 0.900 ;
        RECT 1.645 0.425 1.815 0.730 ;
        RECT 0.965 0.255 1.815 0.425 ;
        RECT 1.985 0.085 2.315 0.560 ;
        RECT 2.485 0.445 2.655 0.730 ;
        RECT 3.155 0.615 3.420 1.410 ;
        RECT 3.590 0.860 3.760 1.750 ;
        RECT 3.970 1.955 4.140 2.285 ;
        RECT 4.335 2.125 4.610 2.455 ;
        RECT 3.970 1.625 4.270 1.955 ;
        RECT 3.930 1.200 4.260 1.415 ;
        RECT 4.440 1.200 4.610 2.125 ;
        RECT 4.780 1.540 4.950 2.625 ;
        RECT 5.120 1.880 5.290 2.735 ;
        RECT 5.510 2.050 5.840 2.905 ;
        RECT 6.200 2.520 6.530 3.245 ;
        RECT 5.120 1.710 5.820 1.880 ;
        RECT 4.780 1.370 5.480 1.540 ;
        RECT 3.930 1.030 5.000 1.200 ;
        RECT 5.170 1.150 5.480 1.370 ;
        RECT 5.650 1.400 5.820 1.710 ;
        RECT 6.050 1.860 6.380 2.240 ;
        RECT 6.760 1.860 7.010 2.700 ;
        RECT 7.210 2.030 7.540 3.245 ;
        RECT 6.050 1.690 7.735 1.860 ;
        RECT 6.050 1.570 6.380 1.690 ;
        RECT 6.875 1.400 7.205 1.520 ;
        RECT 5.650 1.230 7.205 1.400 ;
        RECT 3.590 0.690 4.660 0.860 ;
        RECT 3.590 0.445 3.760 0.690 ;
        RECT 2.485 0.275 3.760 0.445 ;
        RECT 4.070 0.085 4.320 0.520 ;
        RECT 4.490 0.425 4.660 0.690 ;
        RECT 4.830 0.595 5.000 1.030 ;
        RECT 5.650 0.980 5.820 1.230 ;
        RECT 6.875 1.190 7.205 1.230 ;
        RECT 7.375 1.350 7.735 1.690 ;
        RECT 5.220 0.730 5.820 0.980 ;
        RECT 5.565 0.425 5.895 0.510 ;
        RECT 4.490 0.255 5.895 0.425 ;
        RECT 6.230 0.085 6.560 1.060 ;
        RECT 7.375 1.020 7.545 1.350 ;
        RECT 6.790 0.850 7.545 1.020 ;
        RECT 6.790 0.350 7.040 0.850 ;
        RECT 7.220 0.085 7.535 0.680 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__dfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.505 1.780 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.725 2.050 2.055 2.380 ;
        RECT 1.885 1.480 2.055 2.050 ;
        RECT 1.885 1.150 2.275 1.480 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.145 1.665 1.240 ;
        RECT 7.260 1.170 8.635 1.240 ;
        RECT 0.005 1.055 3.445 1.145 ;
        RECT 5.330 1.055 8.635 1.170 ;
        RECT 0.005 0.245 8.635 1.055 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 7.745 2.030 8.105 2.980 ;
        RECT 7.935 1.130 8.105 2.030 ;
        RECT 7.765 0.350 8.105 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.645 2.290 0.815 3.245 ;
        RECT 1.015 2.795 1.345 2.980 ;
        RECT 1.575 2.965 1.935 3.245 ;
        RECT 3.710 2.965 4.100 3.245 ;
        RECT 2.105 2.795 3.540 2.925 ;
        RECT 4.820 2.905 5.875 3.075 ;
        RECT 4.820 2.795 4.990 2.905 ;
        RECT 1.015 2.755 4.990 2.795 ;
        RECT 1.015 2.625 2.275 2.755 ;
        RECT 3.370 2.625 4.990 2.755 ;
        RECT 0.115 1.950 0.845 2.120 ;
        RECT 0.675 1.550 0.845 1.950 ;
        RECT 1.015 1.720 1.475 2.625 ;
        RECT 2.225 1.820 2.555 2.455 ;
        RECT 2.755 2.425 2.955 2.585 ;
        RECT 2.755 2.255 4.135 2.425 ;
        RECT 2.755 2.125 2.955 2.255 ;
        RECT 0.675 1.130 1.135 1.550 ;
        RECT 0.115 0.960 1.135 1.130 ;
        RECT 0.115 0.350 0.365 0.960 ;
        RECT 0.545 0.085 0.795 0.790 ;
        RECT 0.965 0.425 1.135 0.960 ;
        RECT 1.305 1.350 1.715 1.720 ;
        RECT 2.225 1.650 2.615 1.820 ;
        RECT 1.305 0.595 1.475 1.350 ;
        RECT 2.445 1.320 2.615 1.650 ;
        RECT 2.785 1.660 2.955 2.125 ;
        RECT 3.140 1.830 3.540 2.085 ;
        RECT 2.785 1.490 3.200 1.660 ;
        RECT 2.445 1.150 2.860 1.320 ;
        RECT 1.645 0.810 2.520 0.980 ;
        RECT 1.645 0.425 1.815 0.810 ;
        RECT 0.965 0.255 1.815 0.425 ;
        RECT 1.985 0.085 2.180 0.640 ;
        RECT 2.350 0.425 2.520 0.810 ;
        RECT 2.690 0.595 2.860 1.150 ;
        RECT 3.030 0.945 3.200 1.490 ;
        RECT 3.370 1.455 3.540 1.830 ;
        RECT 3.965 1.955 4.135 2.255 ;
        RECT 4.305 2.125 4.650 2.455 ;
        RECT 3.965 1.625 4.310 1.955 ;
        RECT 3.370 1.285 3.755 1.455 ;
        RECT 4.480 1.415 4.650 2.125 ;
        RECT 3.030 0.615 3.415 0.945 ;
        RECT 3.585 0.860 3.755 1.285 ;
        RECT 3.925 1.200 4.650 1.415 ;
        RECT 4.820 1.540 4.990 2.625 ;
        RECT 5.160 1.880 5.330 2.735 ;
        RECT 5.545 2.050 5.875 2.905 ;
        RECT 6.235 2.520 6.565 3.245 ;
        RECT 5.160 1.710 5.755 1.880 ;
        RECT 4.820 1.370 5.415 1.540 ;
        RECT 3.925 1.030 4.915 1.200 ;
        RECT 5.085 1.150 5.415 1.370 ;
        RECT 5.585 1.400 5.755 1.710 ;
        RECT 6.085 1.860 6.415 2.240 ;
        RECT 6.790 1.860 7.040 2.860 ;
        RECT 7.240 2.030 7.570 3.245 ;
        RECT 6.085 1.690 7.765 1.860 ;
        RECT 8.275 1.820 8.525 3.245 ;
        RECT 6.085 1.570 6.415 1.690 ;
        RECT 6.910 1.400 7.240 1.520 ;
        RECT 5.585 1.230 7.240 1.400 ;
        RECT 4.745 0.945 4.915 1.030 ;
        RECT 5.585 0.945 5.755 1.230 ;
        RECT 6.910 1.190 7.240 1.230 ;
        RECT 7.425 1.350 7.765 1.690 ;
        RECT 3.585 0.690 4.575 0.860 ;
        RECT 3.585 0.425 3.755 0.690 ;
        RECT 2.350 0.255 3.755 0.425 ;
        RECT 3.985 0.085 4.235 0.520 ;
        RECT 4.405 0.425 4.575 0.690 ;
        RECT 4.745 0.595 5.075 0.945 ;
        RECT 5.245 0.695 5.755 0.945 ;
        RECT 5.560 0.425 5.890 0.510 ;
        RECT 4.405 0.255 5.890 0.425 ;
        RECT 6.225 0.085 6.555 1.060 ;
        RECT 7.425 1.020 7.595 1.350 ;
        RECT 6.785 0.850 7.595 1.020 ;
        RECT 6.785 0.350 7.115 0.850 ;
        RECT 7.300 0.085 7.595 0.680 ;
        RECT 8.275 0.085 8.525 1.130 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__dfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.505 1.780 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.785 2.025 2.115 2.355 ;
        RECT 1.945 1.780 2.115 2.025 ;
        RECT 1.945 1.125 2.305 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.145 1.665 1.240 ;
        RECT 6.780 1.170 9.570 1.240 ;
        RECT 0.005 1.060 3.580 1.145 ;
        RECT 4.775 1.060 9.570 1.170 ;
        RECT 0.005 0.245 9.570 1.060 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.970 8.135 2.980 ;
        RECT 8.705 1.970 9.035 2.980 ;
        RECT 7.805 1.800 9.035 1.970 ;
        RECT 8.865 1.130 9.035 1.800 ;
        RECT 7.820 0.960 9.035 1.130 ;
        RECT 7.820 0.350 8.150 0.960 ;
        RECT 8.700 0.350 9.035 0.960 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.645 2.290 0.815 3.245 ;
        RECT 1.015 2.695 1.475 2.980 ;
        RECT 1.655 2.865 1.825 3.245 ;
        RECT 1.995 2.905 3.375 3.075 ;
        RECT 3.715 2.930 4.045 3.245 ;
        RECT 1.995 2.695 2.165 2.905 ;
        RECT 3.205 2.760 3.375 2.905 ;
        RECT 4.215 2.905 5.955 3.075 ;
        RECT 4.215 2.760 4.385 2.905 ;
        RECT 1.015 2.525 2.165 2.695 ;
        RECT 0.115 1.950 0.845 2.120 ;
        RECT 0.675 1.550 0.845 1.950 ;
        RECT 1.015 1.820 1.475 2.525 ;
        RECT 2.335 2.120 2.505 2.735 ;
        RECT 2.705 2.485 3.035 2.735 ;
        RECT 3.205 2.590 4.385 2.760 ;
        RECT 2.815 2.420 3.035 2.485 ;
        RECT 2.815 2.250 4.385 2.420 ;
        RECT 2.335 1.950 2.645 2.120 ;
        RECT 1.305 1.550 1.475 1.820 ;
        RECT 0.675 1.130 1.135 1.550 ;
        RECT 0.115 0.960 1.135 1.130 ;
        RECT 0.115 0.350 0.445 0.960 ;
        RECT 0.625 0.085 0.795 0.790 ;
        RECT 0.965 0.425 1.135 0.960 ;
        RECT 1.305 1.220 1.765 1.550 ;
        RECT 2.475 1.240 2.645 1.950 ;
        RECT 2.815 1.580 2.985 2.250 ;
        RECT 3.155 1.750 3.875 2.080 ;
        RECT 2.815 1.410 3.345 1.580 ;
        RECT 1.305 0.595 1.475 1.220 ;
        RECT 2.475 1.070 2.995 1.240 ;
        RECT 1.645 0.730 2.655 0.900 ;
        RECT 1.645 0.425 1.815 0.730 ;
        RECT 0.965 0.255 1.815 0.425 ;
        RECT 1.985 0.085 2.315 0.560 ;
        RECT 2.485 0.425 2.655 0.730 ;
        RECT 2.825 0.595 2.995 1.070 ;
        RECT 3.175 0.950 3.345 1.410 ;
        RECT 3.175 0.620 3.535 0.950 ;
        RECT 3.705 0.860 3.875 1.750 ;
        RECT 4.055 1.630 4.385 2.250 ;
        RECT 4.555 1.370 4.725 2.735 ;
        RECT 4.895 1.540 5.065 2.905 ;
        RECT 5.235 1.880 5.405 2.735 ;
        RECT 5.625 2.050 5.955 2.905 ;
        RECT 6.315 2.450 6.650 3.245 ;
        RECT 6.820 1.890 7.150 2.980 ;
        RECT 7.355 2.060 7.605 3.245 ;
        RECT 8.335 2.140 8.505 3.245 ;
        RECT 5.235 1.710 5.860 1.880 ;
        RECT 6.290 1.810 7.470 1.890 ;
        RECT 9.235 1.820 9.485 3.245 ;
        RECT 4.895 1.370 5.520 1.540 ;
        RECT 4.045 1.200 4.725 1.370 ;
        RECT 4.045 1.030 5.020 1.200 ;
        RECT 5.190 1.150 5.520 1.370 ;
        RECT 5.690 1.310 5.860 1.710 ;
        RECT 6.130 1.720 7.470 1.810 ;
        RECT 6.130 1.480 6.460 1.720 ;
        RECT 7.300 1.630 7.470 1.720 ;
        RECT 6.800 1.390 7.130 1.550 ;
        RECT 6.630 1.310 7.130 1.390 ;
        RECT 5.690 1.220 7.130 1.310 ;
        RECT 7.300 1.300 8.665 1.630 ;
        RECT 4.850 0.950 5.020 1.030 ;
        RECT 5.690 1.140 6.800 1.220 ;
        RECT 5.690 0.970 5.860 1.140 ;
        RECT 7.300 1.050 7.470 1.300 ;
        RECT 6.970 0.970 7.470 1.050 ;
        RECT 3.705 0.690 4.680 0.860 ;
        RECT 3.705 0.425 3.875 0.690 ;
        RECT 2.485 0.255 3.875 0.425 ;
        RECT 4.090 0.085 4.340 0.520 ;
        RECT 4.510 0.425 4.680 0.690 ;
        RECT 4.850 0.595 5.180 0.950 ;
        RECT 5.350 0.720 5.860 0.970 ;
        RECT 5.665 0.425 5.995 0.510 ;
        RECT 4.510 0.255 5.995 0.425 ;
        RECT 6.410 0.085 6.660 0.970 ;
        RECT 6.890 0.880 7.470 0.970 ;
        RECT 6.890 0.350 7.140 0.880 ;
        RECT 7.320 0.085 7.650 0.710 ;
        RECT 8.330 0.085 8.500 0.790 ;
        RECT 9.210 0.085 9.460 1.130 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
  END
END sky130_fd_sc_hs__dfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hs__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641700 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.265 0.865 3.065 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 0.955 1.380 ;
        RECT 0.000 0.000 0.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.150 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.960 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.960 3.415 ;
        RECT 0.000 -0.085 0.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
  END
END sky130_fd_sc_hs__diode_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.459000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.475 5.155 1.805 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.470 1.335 1.800 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.880 1.395 4.825 1.495 ;
        RECT 2.880 1.240 5.725 1.395 ;
        RECT 0.005 1.170 0.950 1.240 ;
        RECT 2.880 1.170 6.715 1.240 ;
        RECT 0.005 0.245 6.715 1.170 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.785 6.910 3.520 ;
        RECT -0.190 1.660 2.670 1.785 ;
        RECT 5.035 1.660 6.910 1.785 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 6.205 1.550 6.605 2.980 ;
        RECT 6.275 0.350 6.605 1.550 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.095 1.820 0.445 2.980 ;
        RECT 0.615 2.310 0.945 3.245 ;
        RECT 1.385 2.550 2.285 2.880 ;
        RECT 2.835 2.730 3.165 3.245 ;
        RECT 3.945 2.560 4.260 2.825 ;
        RECT 1.385 2.140 1.555 2.550 ;
        RECT 3.030 2.390 4.260 2.560 ;
        RECT 3.030 2.380 3.200 2.390 ;
        RECT 0.615 1.970 1.555 2.140 ;
        RECT 1.725 2.050 3.200 2.380 ;
        RECT 3.370 2.050 3.775 2.220 ;
        RECT 0.095 1.130 0.265 1.820 ;
        RECT 0.615 1.630 0.785 1.970 ;
        RECT 0.435 1.300 0.785 1.630 ;
        RECT 0.615 1.130 1.555 1.300 ;
        RECT 1.725 1.150 1.995 2.050 ;
        RECT 2.205 1.330 2.535 1.840 ;
        RECT 3.030 1.830 3.200 2.050 ;
        RECT 3.030 1.500 3.435 1.830 ;
        RECT 3.605 1.330 3.775 2.050 ;
        RECT 2.205 1.160 3.775 1.330 ;
        RECT 0.095 0.960 0.445 1.130 ;
        RECT 1.385 0.980 1.555 1.130 ;
        RECT 0.095 0.790 1.215 0.960 ;
        RECT 0.095 0.350 0.445 0.790 ;
        RECT 0.625 0.085 0.875 0.620 ;
        RECT 1.045 0.425 1.215 0.790 ;
        RECT 1.385 0.650 2.260 0.980 ;
        RECT 2.750 0.685 3.295 0.935 ;
        RECT 2.625 0.425 2.955 0.510 ;
        RECT 1.045 0.255 2.955 0.425 ;
        RECT 3.125 0.085 3.295 0.685 ;
        RECT 3.465 0.605 3.775 1.160 ;
        RECT 3.945 1.945 4.260 2.390 ;
        RECT 4.430 1.975 4.760 3.245 ;
        RECT 4.930 2.145 5.260 2.825 ;
        RECT 4.930 1.975 5.535 2.145 ;
        RECT 3.945 1.055 4.205 1.945 ;
        RECT 5.365 1.630 5.535 1.975 ;
        RECT 5.705 1.945 6.035 3.245 ;
        RECT 4.385 0.085 4.715 1.305 ;
        RECT 5.365 1.300 6.035 1.630 ;
        RECT 5.365 1.285 5.615 1.300 ;
        RECT 5.285 0.605 5.615 1.285 ;
        RECT 5.845 0.085 6.095 1.130 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__dlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlclkp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 4.550 1.445 5.220 1.780 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.450 1.335 1.780 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.200 1.465 4.145 1.495 ;
        RECT 3.200 1.330 5.995 1.465 ;
        RECT 3.200 1.245 7.675 1.330 ;
        RECT 0.005 1.140 0.950 1.240 ;
        RECT 2.415 1.140 7.675 1.245 ;
        RECT 0.005 0.245 7.675 1.140 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.780 7.870 3.520 ;
        RECT -0.190 1.660 1.160 1.780 ;
        RECT 4.355 1.755 7.870 1.780 ;
        RECT 6.205 1.660 7.870 1.755 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 6.805 0.440 7.135 2.980 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.095 1.820 0.445 2.980 ;
        RECT 0.685 2.290 1.075 3.245 ;
        RECT 1.535 2.550 2.405 2.880 ;
        RECT 2.945 2.650 3.485 3.245 ;
        RECT 1.535 2.120 1.705 2.550 ;
        RECT 2.225 2.220 2.555 2.380 ;
        RECT 0.615 1.950 1.705 2.120 ;
        RECT 1.875 2.050 3.325 2.220 ;
        RECT 0.095 0.940 0.265 1.820 ;
        RECT 0.615 1.550 0.785 1.950 ;
        RECT 0.435 1.280 0.785 1.550 ;
        RECT 1.875 1.450 2.045 2.050 ;
        RECT 3.155 1.885 3.325 2.050 ;
        RECT 3.655 2.100 3.985 2.980 ;
        RECT 0.435 1.110 1.560 1.280 ;
        RECT 1.730 1.120 2.045 1.450 ;
        RECT 2.255 1.385 2.585 1.840 ;
        RECT 3.155 1.555 3.485 1.885 ;
        RECT 3.655 1.385 3.825 2.100 ;
        RECT 4.210 2.075 4.545 2.955 ;
        RECT 4.715 2.075 5.045 3.245 ;
        RECT 4.210 1.885 4.380 2.075 ;
        RECT 5.215 1.950 5.560 2.955 ;
        RECT 5.730 1.950 6.635 3.245 ;
        RECT 3.995 1.555 4.380 1.885 ;
        RECT 2.255 1.215 4.035 1.385 ;
        RECT 1.390 0.950 1.560 1.110 ;
        RECT 0.095 0.770 1.220 0.940 ;
        RECT 0.095 0.350 0.365 0.770 ;
        RECT 0.545 0.085 0.880 0.600 ;
        RECT 1.050 0.425 1.220 0.770 ;
        RECT 1.390 0.620 2.245 0.950 ;
        RECT 2.920 0.755 3.535 1.005 ;
        RECT 2.830 0.425 3.160 0.585 ;
        RECT 1.050 0.255 3.160 0.425 ;
        RECT 3.340 0.085 3.535 0.755 ;
        RECT 3.705 0.605 4.035 1.215 ;
        RECT 4.210 1.275 4.380 1.555 ;
        RECT 5.390 1.610 5.560 1.950 ;
        RECT 7.315 1.820 7.565 3.245 ;
        RECT 4.210 0.575 4.595 1.275 ;
        RECT 4.765 0.085 5.095 1.275 ;
        RECT 5.390 0.940 6.305 1.610 ;
        RECT 5.555 0.575 5.885 0.940 ;
        RECT 6.305 0.085 6.635 0.770 ;
        RECT 7.315 0.085 7.565 1.220 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__dlclkp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlclkp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.516000 ;
    PORT
      LAYER li1 ;
        RECT 4.400 1.360 5.070 1.780 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.530 1.430 1.800 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.715 1.495 4.265 1.720 ;
        RECT 2.425 1.240 4.265 1.495 ;
        RECT 0.005 1.170 0.950 1.240 ;
        RECT 2.425 1.170 8.635 1.240 ;
        RECT 0.005 0.245 8.635 1.170 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.930 8.830 3.520 ;
        RECT -0.190 1.705 3.205 1.930 ;
        RECT -0.190 1.660 2.215 1.705 ;
        RECT 4.475 1.660 8.830 1.930 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.103200 ;
    PORT
      LAYER li1 ;
        RECT 6.795 1.720 7.125 2.980 ;
        RECT 7.745 1.780 7.995 2.980 ;
        RECT 7.745 1.720 8.515 1.780 ;
        RECT 6.795 1.550 8.515 1.720 ;
        RECT 7.805 1.380 8.015 1.550 ;
        RECT 6.835 1.210 8.015 1.380 ;
        RECT 6.835 0.350 7.165 1.210 ;
        RECT 7.765 0.350 8.015 1.210 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.115 1.820 0.540 2.980 ;
        RECT 0.785 2.310 1.160 3.245 ;
        RECT 3.110 2.860 3.440 3.245 ;
        RECT 1.435 2.520 2.485 2.850 ;
        RECT 4.205 2.690 4.535 2.970 ;
        RECT 3.305 2.520 4.535 2.690 ;
        RECT 1.435 2.140 1.605 2.520 ;
        RECT 3.305 2.350 3.475 2.520 ;
        RECT 0.710 1.970 1.605 2.140 ;
        RECT 1.775 2.050 3.475 2.350 ;
        RECT 3.645 2.180 3.995 2.350 ;
        RECT 0.115 1.020 0.365 1.820 ;
        RECT 0.710 1.550 0.880 1.970 ;
        RECT 0.535 1.360 0.880 1.550 ;
        RECT 0.535 1.190 1.605 1.360 ;
        RECT 0.115 0.850 1.265 1.020 ;
        RECT 0.115 0.350 0.365 0.850 ;
        RECT 0.550 0.085 0.925 0.680 ;
        RECT 1.095 0.425 1.265 0.850 ;
        RECT 1.435 0.980 1.605 1.190 ;
        RECT 1.775 1.150 2.065 2.050 ;
        RECT 3.305 1.960 3.475 2.050 ;
        RECT 2.305 1.530 2.635 1.805 ;
        RECT 3.305 1.700 3.655 1.960 ;
        RECT 3.825 1.610 3.995 2.180 ;
        RECT 4.205 2.090 4.535 2.520 ;
        RECT 4.740 2.090 5.070 3.245 ;
        RECT 5.240 1.990 5.570 2.980 ;
        RECT 5.740 2.160 6.625 3.245 ;
        RECT 5.240 1.820 6.350 1.990 ;
        RECT 7.295 1.890 7.545 3.245 ;
        RECT 8.195 1.950 8.525 3.245 ;
        RECT 3.825 1.530 4.155 1.610 ;
        RECT 2.305 1.360 4.155 1.530 ;
        RECT 5.260 1.300 5.805 1.630 ;
        RECT 5.260 1.190 5.430 1.300 ;
        RECT 2.815 1.020 5.430 1.190 ;
        RECT 5.975 1.130 6.350 1.820 ;
        RECT 1.435 0.650 2.330 0.980 ;
        RECT 2.815 0.425 3.145 1.020 ;
        RECT 1.095 0.255 3.145 0.425 ;
        RECT 3.315 0.085 3.645 0.850 ;
        RECT 4.280 0.515 4.610 0.850 ;
        RECT 3.815 0.255 4.610 0.515 ;
        RECT 4.780 0.085 5.110 0.850 ;
        RECT 5.600 0.670 6.350 1.130 ;
        RECT 5.600 0.350 5.975 0.670 ;
        RECT 6.160 0.085 6.655 0.500 ;
        RECT 7.335 0.085 7.585 1.040 ;
        RECT 8.195 0.085 8.525 1.040 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__dlclkp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.260 0.835 1.900 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.260 1.335 1.900 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 5.875 1.180 6.180 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 1.140 2.680 1.240 ;
        RECT 5.100 1.140 8.615 1.240 ;
        RECT 0.010 0.245 8.615 1.140 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
        RECT 1.535 1.560 7.080 1.660 ;
        RECT 5.025 1.530 7.080 1.560 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.535700 ;
    PORT
      LAYER li1 ;
        RECT 6.690 1.720 7.115 2.850 ;
        RECT 6.945 1.050 7.115 1.720 ;
        RECT 6.565 0.350 7.115 1.050 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 8.195 1.820 8.530 2.980 ;
        RECT 8.360 1.130 8.530 1.820 ;
        RECT 8.245 0.350 8.530 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.095 2.240 0.365 2.980 ;
        RECT 0.565 2.410 0.895 3.245 ;
        RECT 2.505 2.900 2.835 3.245 ;
        RECT 3.120 2.905 4.290 3.075 ;
        RECT 1.065 2.730 2.015 2.900 ;
        RECT 1.065 2.240 1.235 2.730 ;
        RECT 1.845 2.560 2.910 2.730 ;
        RECT 0.095 2.070 1.235 2.240 ;
        RECT 1.405 2.390 1.675 2.560 ;
        RECT 1.405 2.220 2.555 2.390 ;
        RECT 1.405 2.100 1.675 2.220 ;
        RECT 0.095 1.090 0.265 2.070 ;
        RECT 1.505 1.090 1.675 2.100 ;
        RECT 0.095 0.540 0.450 1.090 ;
        RECT 0.630 0.085 0.960 1.090 ;
        RECT 1.130 0.350 1.675 1.090 ;
        RECT 1.845 1.720 2.215 2.050 ;
        RECT 1.845 0.960 2.015 1.720 ;
        RECT 2.385 1.550 2.555 2.220 ;
        RECT 2.185 1.300 2.555 1.550 ;
        RECT 2.740 1.800 2.910 2.560 ;
        RECT 3.120 2.140 3.290 2.905 ;
        RECT 3.460 2.405 3.790 2.735 ;
        RECT 3.120 1.970 3.450 2.140 ;
        RECT 2.740 1.470 3.070 1.800 ;
        RECT 3.280 1.450 3.450 1.970 ;
        RECT 3.620 1.790 3.790 2.405 ;
        RECT 3.960 2.050 4.290 2.905 ;
        RECT 4.680 2.520 5.445 3.245 ;
        RECT 5.615 2.290 5.945 2.850 ;
        RECT 4.530 1.960 5.945 2.290 ;
        RECT 6.115 2.060 6.445 3.245 ;
        RECT 5.290 1.890 5.945 1.960 ;
        RECT 3.620 1.620 4.725 1.790 ;
        RECT 4.375 1.550 4.725 1.620 ;
        RECT 5.290 1.720 6.520 1.890 ;
        RECT 3.280 1.300 3.610 1.450 ;
        RECT 2.185 1.130 3.610 1.300 ;
        RECT 3.280 1.120 3.610 1.130 ;
        RECT 1.845 0.950 2.175 0.960 ;
        RECT 3.875 0.950 4.205 1.450 ;
        RECT 1.845 0.780 4.205 0.950 ;
        RECT 4.375 1.220 5.120 1.550 ;
        RECT 1.845 0.350 2.175 0.780 ;
        RECT 4.375 0.610 4.545 1.220 ;
        RECT 5.290 1.050 5.460 1.720 ;
        RECT 6.350 1.550 6.520 1.720 ;
        RECT 7.285 1.630 7.535 2.780 ;
        RECT 7.745 1.820 8.010 3.245 ;
        RECT 6.350 1.220 6.775 1.550 ;
        RECT 7.285 1.300 8.190 1.630 ;
        RECT 2.345 0.085 2.915 0.600 ;
        RECT 3.405 0.360 4.545 0.610 ;
        RECT 4.730 0.085 4.980 1.030 ;
        RECT 5.210 0.350 5.460 1.050 ;
        RECT 6.030 0.085 6.360 1.010 ;
        RECT 7.285 0.540 7.560 1.300 ;
        RECT 7.745 0.085 8.075 1.130 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__dlrbn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.260 0.805 1.930 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.260 1.285 1.930 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 5.570 1.180 6.115 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 2.630 1.240 ;
        RECT 0.005 0.920 3.730 1.140 ;
        RECT 4.765 0.920 9.115 1.240 ;
        RECT 0.005 0.245 9.115 0.920 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
        RECT 1.455 1.560 2.295 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 6.260 1.820 6.590 2.070 ;
        RECT 6.285 1.130 6.455 1.820 ;
        RECT 6.285 0.770 6.615 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.572800 ;
    PORT
      LAYER li1 ;
        RECT 8.225 1.820 8.575 2.980 ;
        RECT 8.405 1.050 8.575 1.820 ;
        RECT 8.205 0.880 8.575 1.050 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.085 2.270 0.445 2.980 ;
        RECT 0.645 2.440 0.815 3.245 ;
        RECT 2.425 2.820 2.755 3.245 ;
        RECT 3.010 2.905 4.165 3.075 ;
        RECT 0.985 2.650 1.965 2.820 ;
        RECT 0.985 2.270 1.155 2.650 ;
        RECT 1.795 2.480 2.830 2.650 ;
        RECT 0.085 2.100 1.155 2.270 ;
        RECT 1.325 2.310 1.625 2.480 ;
        RECT 1.325 2.140 2.475 2.310 ;
        RECT 1.325 2.100 1.625 2.140 ;
        RECT 0.085 1.090 0.255 2.100 ;
        RECT 1.455 1.090 1.625 2.100 ;
        RECT 0.085 0.540 0.445 1.090 ;
        RECT 0.625 0.085 0.955 1.090 ;
        RECT 1.125 0.350 1.625 1.090 ;
        RECT 1.795 1.720 2.135 1.970 ;
        RECT 1.795 0.960 1.965 1.720 ;
        RECT 2.305 1.550 2.475 2.140 ;
        RECT 2.135 1.300 2.475 1.550 ;
        RECT 2.660 1.800 2.830 2.480 ;
        RECT 3.010 2.140 3.180 2.905 ;
        RECT 3.350 2.405 3.665 2.735 ;
        RECT 3.010 1.970 3.325 2.140 ;
        RECT 2.660 1.470 2.985 1.800 ;
        RECT 3.155 1.450 3.325 1.970 ;
        RECT 3.495 1.880 3.665 2.405 ;
        RECT 3.835 2.050 4.165 2.905 ;
        RECT 4.525 2.650 5.140 3.245 ;
        RECT 5.310 2.410 5.640 2.980 ;
        RECT 5.810 2.580 6.140 3.245 ;
        RECT 6.710 2.580 7.040 3.245 ;
        RECT 5.310 2.350 6.955 2.410 ;
        RECT 4.375 2.240 6.955 2.350 ;
        RECT 4.375 2.050 5.640 2.240 ;
        RECT 3.495 1.710 5.060 1.880 ;
        RECT 3.155 1.300 3.530 1.450 ;
        RECT 2.135 1.130 3.530 1.300 ;
        RECT 3.155 1.120 3.530 1.130 ;
        RECT 3.715 1.225 4.130 1.540 ;
        RECT 1.795 0.950 2.125 0.960 ;
        RECT 3.715 0.950 3.885 1.225 ;
        RECT 4.300 1.055 4.470 1.710 ;
        RECT 4.735 1.350 5.060 1.710 ;
        RECT 5.230 1.820 5.640 2.050 ;
        RECT 5.230 1.130 5.400 1.820 ;
        RECT 6.785 1.650 6.955 2.240 ;
        RECT 6.625 1.320 6.955 1.650 ;
        RECT 7.215 1.550 7.545 2.860 ;
        RECT 7.775 1.820 8.025 3.245 ;
        RECT 8.755 1.820 9.005 3.245 ;
        RECT 1.795 0.780 3.885 0.950 ;
        RECT 4.055 0.885 4.470 1.055 ;
        RECT 1.795 0.350 2.125 0.780 ;
        RECT 4.055 0.610 4.225 0.885 ;
        RECT 2.295 0.085 2.835 0.600 ;
        RECT 3.325 0.360 4.225 0.610 ;
        RECT 4.395 0.085 4.645 0.715 ;
        RECT 4.875 0.350 5.400 1.130 ;
        RECT 7.215 1.220 8.230 1.550 ;
        RECT 5.695 0.085 6.025 1.010 ;
        RECT 6.785 0.085 7.045 1.050 ;
        RECT 7.215 0.350 7.545 1.220 ;
        RECT 7.775 0.085 8.035 1.050 ;
        RECT 8.745 0.085 9.005 1.130 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__dlrbn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.450 0.805 1.780 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.450 1.305 1.780 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 5.425 1.180 5.795 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.360 1.625 1.390 ;
        RECT 0.005 1.170 2.645 1.360 ;
        RECT 4.690 1.170 8.155 1.240 ;
        RECT 0.005 0.245 8.155 1.170 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 6.200 2.060 6.670 2.980 ;
        RECT 6.500 1.180 6.670 2.060 ;
        RECT 6.130 1.010 6.670 1.180 ;
        RECT 6.130 0.350 6.460 1.010 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.604200 ;
    PORT
      LAYER li1 ;
        RECT 7.715 1.820 8.055 2.980 ;
        RECT 7.885 1.040 8.055 1.820 ;
        RECT 7.710 0.350 8.055 1.040 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.095 2.560 0.445 2.850 ;
        RECT 0.650 2.730 0.980 3.245 ;
        RECT 2.350 2.730 2.685 3.245 ;
        RECT 2.855 2.905 4.015 3.075 ;
        RECT 0.095 2.390 2.675 2.560 ;
        RECT 0.095 1.970 0.445 2.390 ;
        RECT 1.185 1.970 1.645 2.220 ;
        RECT 0.095 1.280 0.265 1.970 ;
        RECT 1.475 1.750 1.645 1.970 ;
        RECT 1.815 1.940 2.215 2.220 ;
        RECT 1.475 1.420 1.875 1.750 ;
        RECT 1.475 1.280 1.645 1.420 ;
        RECT 0.095 0.690 0.445 1.280 ;
        RECT 0.625 0.085 0.955 1.280 ;
        RECT 1.185 0.750 1.645 1.280 ;
        RECT 2.045 1.300 2.215 1.940 ;
        RECT 2.505 1.800 2.675 2.390 ;
        RECT 2.855 2.140 3.025 2.905 ;
        RECT 3.195 2.405 3.515 2.735 ;
        RECT 2.855 1.970 3.175 2.140 ;
        RECT 2.505 1.470 2.835 1.800 ;
        RECT 3.005 1.480 3.175 1.970 ;
        RECT 3.345 1.820 3.515 2.405 ;
        RECT 3.685 2.050 4.015 2.905 ;
        RECT 4.405 2.650 5.080 3.245 ;
        RECT 5.250 2.320 5.580 2.980 ;
        RECT 4.225 1.990 5.580 2.320 ;
        RECT 5.780 2.060 6.030 3.245 ;
        RECT 5.085 1.890 5.580 1.990 ;
        RECT 3.345 1.650 4.915 1.820 ;
        RECT 3.005 1.300 3.395 1.480 ;
        RECT 2.045 1.250 3.395 1.300 ;
        RECT 1.825 1.130 3.395 1.250 ;
        RECT 1.825 0.920 2.215 1.130 ;
        RECT 3.580 0.960 3.750 1.650 ;
        RECT 4.585 1.350 4.915 1.650 ;
        RECT 5.085 1.720 6.330 1.890 ;
        RECT 5.085 1.130 5.255 1.720 ;
        RECT 6.005 1.350 6.330 1.720 ;
        RECT 6.840 1.650 7.010 2.980 ;
        RECT 7.210 2.100 7.540 3.245 ;
        RECT 1.185 0.580 2.990 0.750 ;
        RECT 3.190 0.710 3.750 0.960 ;
        RECT 1.185 0.500 1.645 0.580 ;
        RECT 2.820 0.510 2.990 0.580 ;
        RECT 2.320 0.085 2.650 0.410 ;
        RECT 2.820 0.255 3.905 0.510 ;
        RECT 4.240 0.085 4.570 1.060 ;
        RECT 4.800 0.350 5.255 1.130 ;
        RECT 6.840 1.320 7.715 1.650 ;
        RECT 5.620 0.085 5.950 1.010 ;
        RECT 6.840 0.840 7.020 1.320 ;
        RECT 6.690 0.350 7.020 0.840 ;
        RECT 7.200 0.085 7.530 0.940 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__dlrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.450 0.805 1.780 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.180 1.285 1.550 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 5.435 1.180 5.785 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.685 1.240 2.630 1.280 ;
        RECT 0.005 1.170 2.630 1.240 ;
        RECT 4.680 1.170 9.115 1.240 ;
        RECT 0.005 0.245 9.115 1.170 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 6.295 1.970 6.465 2.980 ;
        RECT 6.295 1.800 7.075 1.970 ;
        RECT 6.845 1.130 7.075 1.800 ;
        RECT 6.150 0.960 7.075 1.130 ;
        RECT 6.150 0.350 6.480 0.960 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 8.225 1.820 8.585 2.980 ;
        RECT 8.415 1.130 8.585 1.820 ;
        RECT 8.245 0.350 8.585 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.085 2.530 0.445 2.820 ;
        RECT 0.650 2.700 0.980 3.245 ;
        RECT 2.330 2.700 2.695 3.245 ;
        RECT 2.975 2.905 4.035 3.075 ;
        RECT 0.085 2.360 2.805 2.530 ;
        RECT 0.085 1.950 0.445 2.360 ;
        RECT 0.085 1.130 0.255 1.950 ;
        RECT 1.185 1.940 1.625 2.190 ;
        RECT 1.795 1.940 2.205 2.190 ;
        RECT 1.455 1.670 1.625 1.940 ;
        RECT 1.455 1.340 1.865 1.670 ;
        RECT 0.085 0.540 0.445 1.130 ;
        RECT 1.455 1.010 1.625 1.340 ;
        RECT 2.035 1.300 2.205 1.940 ;
        RECT 2.485 1.470 2.805 2.360 ;
        RECT 2.975 1.480 3.145 2.905 ;
        RECT 3.315 1.820 3.485 2.735 ;
        RECT 3.705 2.050 4.035 2.905 ;
        RECT 4.425 2.650 5.065 3.245 ;
        RECT 5.235 2.320 5.565 2.980 ;
        RECT 4.245 1.990 5.565 2.320 ;
        RECT 5.735 2.060 6.065 3.245 ;
        RECT 6.665 2.140 6.995 3.245 ;
        RECT 5.095 1.890 5.565 1.990 ;
        RECT 3.315 1.650 4.925 1.820 ;
        RECT 2.975 1.300 3.385 1.480 ;
        RECT 2.035 1.170 3.385 1.300 ;
        RECT 0.625 0.085 0.955 1.010 ;
        RECT 1.125 0.750 1.625 1.010 ;
        RECT 1.795 1.130 3.385 1.170 ;
        RECT 1.795 0.920 2.205 1.130 ;
        RECT 3.570 0.960 3.740 1.650 ;
        RECT 4.605 1.350 4.925 1.650 ;
        RECT 5.095 1.720 6.125 1.890 ;
        RECT 5.095 1.130 5.265 1.720 ;
        RECT 5.955 1.630 6.125 1.720 ;
        RECT 7.245 1.630 7.555 2.860 ;
        RECT 7.725 1.820 8.055 3.245 ;
        RECT 8.755 1.820 9.005 3.245 ;
        RECT 5.955 1.300 6.650 1.630 ;
        RECT 7.245 1.300 8.245 1.630 ;
        RECT 3.180 0.790 3.740 0.960 ;
        RECT 1.125 0.580 2.980 0.750 ;
        RECT 1.125 0.350 1.625 0.580 ;
        RECT 2.810 0.510 2.980 0.580 ;
        RECT 2.305 0.085 2.640 0.410 ;
        RECT 2.810 0.255 3.895 0.510 ;
        RECT 4.230 0.085 4.560 1.060 ;
        RECT 4.790 0.350 5.265 1.130 ;
        RECT 7.245 1.130 7.555 1.300 ;
        RECT 5.610 0.085 5.940 1.010 ;
        RECT 6.650 0.085 6.980 0.790 ;
        RECT 7.245 0.450 7.575 1.130 ;
        RECT 7.745 0.085 8.075 1.130 ;
        RECT 8.755 0.085 9.005 1.130 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__dlrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.450 0.835 1.780 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.450 1.335 1.780 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.180 6.235 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.280 1.555 1.360 ;
        RECT 0.005 1.140 2.680 1.280 ;
        RECT 0.005 0.920 4.175 1.140 ;
        RECT 5.130 0.920 7.170 1.240 ;
        RECT 0.005 0.245 7.170 0.920 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.600500 ;
    PORT
      LAYER li1 ;
        RECT 6.755 1.820 7.115 2.980 ;
        RECT 6.945 1.130 7.115 1.820 ;
        RECT 6.730 0.350 7.115 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.095 1.950 0.450 2.830 ;
        RECT 0.655 1.950 0.985 3.245 ;
        RECT 2.300 2.860 2.630 3.245 ;
        RECT 1.190 2.690 1.675 2.830 ;
        RECT 1.190 2.520 4.245 2.690 ;
        RECT 4.635 2.530 5.430 3.245 ;
        RECT 1.190 1.950 1.675 2.520 ;
        RECT 0.095 1.250 0.265 1.950 ;
        RECT 1.505 1.670 1.675 1.950 ;
        RECT 1.845 2.010 2.245 2.350 ;
        RECT 3.255 2.180 3.745 2.350 ;
        RECT 1.845 1.840 3.405 2.010 ;
        RECT 1.505 1.340 1.905 1.670 ;
        RECT 1.505 1.250 1.675 1.340 ;
        RECT 0.095 0.750 0.445 1.250 ;
        RECT 1.065 0.920 1.675 1.250 ;
        RECT 2.075 1.170 2.245 1.840 ;
        RECT 1.845 0.920 2.245 1.170 ;
        RECT 2.535 0.750 2.865 1.590 ;
        RECT 3.075 1.520 3.405 1.840 ;
        RECT 3.575 1.860 3.745 2.180 ;
        RECT 3.915 2.030 4.245 2.520 ;
        RECT 5.635 2.360 5.965 2.860 ;
        RECT 4.485 2.030 5.965 2.360 ;
        RECT 6.255 2.060 6.585 3.245 ;
        RECT 5.465 1.890 5.965 2.030 ;
        RECT 3.575 1.690 5.070 1.860 ;
        RECT 4.900 1.630 5.070 1.690 ;
        RECT 5.465 1.720 6.585 1.890 ;
        RECT 3.075 1.190 4.335 1.520 ;
        RECT 4.900 1.300 5.295 1.630 ;
        RECT 4.900 1.020 5.070 1.300 ;
        RECT 5.465 1.130 5.635 1.720 ;
        RECT 6.415 1.650 6.585 1.720 ;
        RECT 6.415 1.320 6.775 1.650 ;
        RECT 0.095 0.580 2.865 0.750 ;
        RECT 3.815 0.850 5.070 1.020 ;
        RECT 0.625 0.085 0.955 0.410 ;
        RECT 2.355 0.085 3.200 0.410 ;
        RECT 3.815 0.350 4.145 0.850 ;
        RECT 4.670 0.085 5.010 0.680 ;
        RECT 5.240 0.350 5.635 1.130 ;
        RECT 6.140 0.085 6.470 1.010 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__dlrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.450 0.835 1.780 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.450 1.335 1.780 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.180 6.305 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.280 1.595 1.360 ;
        RECT 0.005 1.140 2.705 1.280 ;
        RECT 0.005 0.920 4.255 1.140 ;
        RECT 5.200 0.920 8.145 1.240 ;
        RECT 0.005 0.245 8.145 0.920 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.820 7.535 2.980 ;
        RECT 7.365 1.470 7.535 1.820 ;
        RECT 7.205 0.350 7.535 1.470 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.095 1.950 0.615 2.830 ;
        RECT 0.785 1.950 1.115 3.245 ;
        RECT 2.380 2.860 2.710 3.245 ;
        RECT 1.285 2.690 1.675 2.830 ;
        RECT 1.285 2.520 4.325 2.690 ;
        RECT 4.715 2.630 5.545 3.245 ;
        RECT 1.285 1.950 1.675 2.520 ;
        RECT 0.095 1.250 0.265 1.950 ;
        RECT 1.505 1.670 1.675 1.950 ;
        RECT 1.845 2.010 2.245 2.350 ;
        RECT 3.335 2.180 3.825 2.350 ;
        RECT 1.845 1.840 3.485 2.010 ;
        RECT 1.505 1.340 1.905 1.670 ;
        RECT 1.505 1.250 1.675 1.340 ;
        RECT 0.095 0.750 0.445 1.250 ;
        RECT 1.135 0.920 1.675 1.250 ;
        RECT 2.075 1.170 2.245 1.840 ;
        RECT 1.845 0.920 2.245 1.170 ;
        RECT 2.615 0.750 2.945 1.590 ;
        RECT 3.155 1.520 3.485 1.840 ;
        RECT 3.655 1.860 3.825 2.180 ;
        RECT 3.995 2.030 4.325 2.520 ;
        RECT 5.715 2.360 6.045 2.980 ;
        RECT 4.565 2.030 6.045 2.360 ;
        RECT 6.320 2.060 6.650 3.245 ;
        RECT 5.545 1.890 6.045 2.030 ;
        RECT 3.655 1.690 5.375 1.860 ;
        RECT 3.155 1.190 4.415 1.520 ;
        RECT 4.970 1.350 5.375 1.690 ;
        RECT 5.545 1.720 6.675 1.890 ;
        RECT 7.705 1.820 8.045 3.245 ;
        RECT 4.970 1.020 5.140 1.350 ;
        RECT 5.545 1.130 5.715 1.720 ;
        RECT 6.505 1.650 6.675 1.720 ;
        RECT 6.505 1.320 6.845 1.650 ;
        RECT 0.095 0.580 2.945 0.750 ;
        RECT 3.895 0.850 5.140 1.020 ;
        RECT 0.625 0.085 0.955 0.410 ;
        RECT 2.380 0.085 3.280 0.410 ;
        RECT 3.895 0.350 4.225 0.850 ;
        RECT 4.750 0.085 5.080 0.680 ;
        RECT 5.310 0.350 5.715 1.130 ;
        RECT 6.130 0.085 7.035 1.010 ;
        RECT 7.705 0.085 8.035 1.130 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__dlrtn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.450 0.805 1.780 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.450 1.290 1.780 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 6.320 1.120 7.555 1.450 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 2.635 1.360 ;
        RECT 7.325 1.140 9.595 1.240 ;
        RECT 0.005 0.920 4.100 1.140 ;
        RECT 5.045 0.920 9.595 1.140 ;
        RECT 0.005 0.245 9.595 0.920 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.198400 ;
    PORT
      LAYER li1 ;
        RECT 7.545 2.130 7.875 2.980 ;
        RECT 8.545 2.130 8.875 2.980 ;
        RECT 7.545 1.970 8.875 2.130 ;
        RECT 7.545 1.960 9.475 1.970 ;
        RECT 8.545 1.800 9.475 1.960 ;
        RECT 9.245 1.130 9.475 1.800 ;
        RECT 7.935 0.960 9.475 1.130 ;
        RECT 7.935 0.360 8.125 0.960 ;
        RECT 8.795 0.800 9.475 0.960 ;
        RECT 8.795 0.360 8.985 0.800 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.085 1.950 0.475 2.830 ;
        RECT 0.645 1.950 0.975 3.245 ;
        RECT 2.255 2.940 2.585 3.245 ;
        RECT 1.145 2.770 1.630 2.830 ;
        RECT 1.145 2.600 4.200 2.770 ;
        RECT 4.590 2.630 5.320 3.245 ;
        RECT 1.145 1.950 1.630 2.600 ;
        RECT 0.085 1.250 0.255 1.950 ;
        RECT 1.460 1.750 1.630 1.950 ;
        RECT 1.800 2.090 2.205 2.430 ;
        RECT 3.180 2.260 3.700 2.430 ;
        RECT 1.800 1.920 3.360 2.090 ;
        RECT 1.460 1.420 1.865 1.750 ;
        RECT 1.460 1.250 1.630 1.420 ;
        RECT 2.035 1.250 2.205 1.920 ;
        RECT 0.085 0.830 0.445 1.250 ;
        RECT 1.135 1.000 1.630 1.250 ;
        RECT 1.800 1.000 2.205 1.250 ;
        RECT 2.490 0.830 2.820 1.670 ;
        RECT 3.030 1.520 3.360 1.920 ;
        RECT 3.530 1.860 3.700 2.260 ;
        RECT 3.870 2.030 4.200 2.600 ;
        RECT 5.490 2.360 5.820 2.960 ;
        RECT 4.440 2.030 5.820 2.360 ;
        RECT 5.990 2.080 6.320 3.245 ;
        RECT 3.530 1.690 5.220 1.860 ;
        RECT 3.030 1.190 4.260 1.520 ;
        RECT 4.815 1.120 5.220 1.690 ;
        RECT 5.490 1.790 5.820 2.030 ;
        RECT 6.490 1.790 6.820 2.960 ;
        RECT 7.045 2.080 7.375 3.245 ;
        RECT 8.045 2.300 8.375 3.245 ;
        RECT 9.045 2.140 9.375 3.245 ;
        RECT 5.490 1.630 7.895 1.790 ;
        RECT 5.490 1.620 9.075 1.630 ;
        RECT 4.815 1.020 4.985 1.120 ;
        RECT 0.085 0.660 2.820 0.830 ;
        RECT 3.740 0.850 4.985 1.020 ;
        RECT 0.625 0.085 0.955 0.490 ;
        RECT 2.310 0.085 3.125 0.490 ;
        RECT 3.740 0.400 4.070 0.850 ;
        RECT 4.595 0.085 4.925 0.680 ;
        RECT 5.155 0.425 5.485 0.950 ;
        RECT 5.665 0.595 5.835 1.620 ;
        RECT 7.725 1.300 9.075 1.620 ;
        RECT 6.015 0.770 7.205 0.950 ;
        RECT 6.015 0.425 6.265 0.770 ;
        RECT 5.155 0.255 6.265 0.425 ;
        RECT 6.445 0.085 6.775 0.600 ;
        RECT 6.945 0.355 7.205 0.770 ;
        RECT 7.435 0.085 7.765 0.950 ;
        RECT 8.295 0.085 8.625 0.790 ;
        RECT 9.155 0.085 9.485 0.630 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
  END
END sky130_fd_sc_hs__dlrtn_4

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.375 1.780 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.930 1.450 1.285 1.780 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 5.435 1.350 5.765 1.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.685 1.240 2.220 1.470 ;
        RECT 0.110 1.140 2.695 1.240 ;
        RECT 0.110 0.920 3.750 1.140 ;
        RECT 4.660 0.920 6.540 1.240 ;
        RECT 0.110 0.245 6.540 0.920 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.780 6.910 3.520 ;
        RECT -0.190 1.660 1.160 1.780 ;
        RECT 2.905 1.660 6.910 1.780 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 6.275 1.820 6.635 2.980 ;
        RECT 6.465 0.840 6.635 1.820 ;
        RECT 6.100 0.350 6.635 0.840 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.115 2.560 0.445 2.980 ;
        RECT 0.615 2.730 0.945 3.245 ;
        RECT 2.330 2.730 2.705 3.245 ;
        RECT 2.905 2.905 4.045 3.075 ;
        RECT 0.115 2.390 2.695 2.560 ;
        RECT 0.115 2.100 0.715 2.390 ;
        RECT 0.545 1.130 0.715 2.100 ;
        RECT 1.150 1.970 1.625 2.220 ;
        RECT 1.795 2.020 2.170 2.220 ;
        RECT 1.455 1.780 1.625 1.970 ;
        RECT 1.455 1.450 1.830 1.780 ;
        RECT 1.455 1.130 1.625 1.450 ;
        RECT 2.000 1.280 2.170 2.020 ;
        RECT 2.525 1.800 2.695 2.390 ;
        RECT 2.905 2.140 3.075 2.905 ;
        RECT 3.245 2.405 3.535 2.735 ;
        RECT 2.905 1.970 3.195 2.140 ;
        RECT 2.525 1.470 2.855 1.800 ;
        RECT 3.025 1.450 3.195 1.970 ;
        RECT 3.365 1.895 3.535 2.405 ;
        RECT 3.715 2.065 4.045 2.905 ;
        RECT 4.435 2.650 5.075 3.245 ;
        RECT 5.245 2.380 5.575 2.980 ;
        RECT 4.305 2.065 5.575 2.380 ;
        RECT 5.095 1.950 5.575 2.065 ;
        RECT 5.745 1.950 6.075 3.245 ;
        RECT 3.365 1.725 4.925 1.895 ;
        RECT 3.025 1.280 3.325 1.450 ;
        RECT 0.220 0.540 0.715 1.130 ;
        RECT 0.885 0.085 1.055 1.130 ;
        RECT 1.235 0.940 1.625 1.130 ;
        RECT 1.795 1.110 3.325 1.280 ;
        RECT 1.235 0.770 3.020 0.940 ;
        RECT 3.495 0.925 3.665 1.725 ;
        RECT 1.235 0.350 1.625 0.770 ;
        RECT 2.295 0.085 2.680 0.600 ;
        RECT 2.850 0.425 3.020 0.770 ;
        RECT 3.190 0.595 3.665 0.925 ;
        RECT 3.835 1.225 4.095 1.555 ;
        RECT 4.665 1.470 4.925 1.725 ;
        RECT 3.835 0.425 4.005 1.225 ;
        RECT 5.095 1.180 5.265 1.950 ;
        RECT 5.975 1.180 6.295 1.550 ;
        RECT 4.770 1.010 6.295 1.180 ;
        RECT 2.850 0.255 4.005 0.425 ;
        RECT 4.210 0.085 4.540 0.810 ;
        RECT 4.770 0.350 5.100 1.010 ;
        RECT 5.590 0.085 5.920 0.840 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__dlrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.515 1.780 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.180 1.285 1.550 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 5.435 1.180 5.840 1.550 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.605 1.240 2.630 1.360 ;
        RECT 0.030 1.140 2.630 1.240 ;
        RECT 0.030 0.955 3.825 1.140 ;
        RECT 4.735 0.955 7.195 1.240 ;
        RECT 0.030 0.245 7.195 0.955 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.567400 ;
    PORT
      LAYER li1 ;
        RECT 6.255 2.060 6.585 2.980 ;
        RECT 6.415 1.970 6.585 2.060 ;
        RECT 6.415 1.800 7.075 1.970 ;
        RECT 6.845 1.130 7.075 1.800 ;
        RECT 6.255 0.960 7.075 1.130 ;
        RECT 6.255 0.350 6.585 0.960 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.115 2.610 0.445 2.820 ;
        RECT 0.650 2.780 0.980 3.245 ;
        RECT 2.280 2.780 2.610 3.245 ;
        RECT 2.890 2.905 4.060 3.075 ;
        RECT 0.115 2.440 2.680 2.610 ;
        RECT 0.115 1.950 0.855 2.440 ;
        RECT 0.685 1.280 0.855 1.950 ;
        RECT 1.185 1.940 1.625 2.270 ;
        RECT 1.825 1.940 2.230 2.270 ;
        RECT 0.140 1.110 0.855 1.280 ;
        RECT 1.455 1.750 1.625 1.940 ;
        RECT 1.455 1.420 1.890 1.750 ;
        RECT 0.140 0.540 0.470 1.110 ;
        RECT 1.455 1.010 1.625 1.420 ;
        RECT 2.060 1.250 2.230 1.940 ;
        RECT 2.510 1.770 2.680 2.440 ;
        RECT 2.890 2.110 3.060 2.905 ;
        RECT 3.230 2.405 3.560 2.735 ;
        RECT 2.890 1.940 3.220 2.110 ;
        RECT 2.510 1.440 2.840 1.770 ;
        RECT 3.050 1.450 3.220 1.940 ;
        RECT 3.390 1.930 3.560 2.405 ;
        RECT 3.730 2.100 4.060 2.905 ;
        RECT 4.450 2.650 5.085 3.245 ;
        RECT 5.255 2.380 5.585 2.980 ;
        RECT 4.300 2.100 5.585 2.380 ;
        RECT 3.390 1.760 4.925 1.930 ;
        RECT 3.050 1.250 3.315 1.450 ;
        RECT 0.650 0.085 0.980 0.940 ;
        RECT 1.150 0.750 1.625 1.010 ;
        RECT 1.795 1.080 3.315 1.250 ;
        RECT 1.795 0.920 2.230 1.080 ;
        RECT 3.485 0.845 3.655 1.760 ;
        RECT 3.825 1.260 4.090 1.590 ;
        RECT 4.660 1.350 4.925 1.760 ;
        RECT 5.095 1.890 5.585 2.100 ;
        RECT 5.755 2.060 6.085 3.245 ;
        RECT 6.755 2.140 7.085 3.245 ;
        RECT 5.095 1.720 6.220 1.890 ;
        RECT 1.150 0.580 2.975 0.750 ;
        RECT 3.205 0.595 3.715 0.845 ;
        RECT 1.150 0.350 1.625 0.580 ;
        RECT 2.805 0.425 2.975 0.580 ;
        RECT 3.920 0.425 4.090 1.260 ;
        RECT 5.095 1.130 5.265 1.720 ;
        RECT 6.050 1.630 6.220 1.720 ;
        RECT 6.050 1.300 6.675 1.630 ;
        RECT 2.305 0.085 2.635 0.410 ;
        RECT 2.805 0.255 4.090 0.425 ;
        RECT 4.285 0.085 4.615 0.845 ;
        RECT 4.845 0.350 5.265 1.130 ;
        RECT 5.755 0.085 6.085 1.010 ;
        RECT 6.755 0.085 7.085 0.790 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__dlrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.515 1.780 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.450 1.290 1.780 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.120 6.595 1.450 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.690 1.310 2.660 1.470 ;
        RECT 0.005 1.140 2.660 1.310 ;
        RECT 6.845 1.140 9.115 1.240 ;
        RECT 0.005 0.920 3.680 1.140 ;
        RECT 4.560 0.920 9.115 1.140 ;
        RECT 0.005 0.245 9.115 0.920 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.780 9.310 3.520 ;
        RECT -0.190 1.660 1.480 1.780 ;
        RECT 2.870 1.660 9.310 1.780 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.164800 ;
    PORT
      LAYER li1 ;
        RECT 7.175 1.970 7.425 2.980 ;
        RECT 8.095 1.970 8.425 2.980 ;
        RECT 7.175 1.800 8.995 1.970 ;
        RECT 8.765 1.130 8.995 1.800 ;
        RECT 7.385 0.880 8.995 1.130 ;
        RECT 7.385 0.365 7.645 0.880 ;
        RECT 8.315 0.365 8.505 0.880 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.115 2.540 0.445 2.830 ;
        RECT 0.650 2.710 0.980 3.245 ;
        RECT 2.335 2.710 2.665 3.245 ;
        RECT 2.845 2.905 3.985 3.075 ;
        RECT 0.115 2.370 2.665 2.540 ;
        RECT 0.115 1.950 0.855 2.370 ;
        RECT 1.185 1.950 1.630 2.200 ;
        RECT 1.800 2.020 2.240 2.200 ;
        RECT 0.685 1.280 0.855 1.950 ;
        RECT 0.115 1.110 0.855 1.280 ;
        RECT 1.460 1.780 1.630 1.950 ;
        RECT 1.460 1.450 1.900 1.780 ;
        RECT 1.460 1.200 1.630 1.450 ;
        RECT 2.070 1.280 2.240 2.020 ;
        RECT 2.495 1.800 2.665 2.370 ;
        RECT 2.845 2.140 3.015 2.905 ;
        RECT 3.185 2.405 3.465 2.735 ;
        RECT 2.845 1.970 3.125 2.140 ;
        RECT 2.495 1.470 2.785 1.800 ;
        RECT 2.955 1.450 3.125 1.970 ;
        RECT 3.295 1.895 3.465 2.405 ;
        RECT 3.655 2.065 3.985 2.905 ;
        RECT 4.345 2.650 4.905 3.245 ;
        RECT 5.110 2.480 5.440 2.700 ;
        RECT 4.195 2.065 5.440 2.480 ;
        RECT 3.295 1.725 5.020 1.895 ;
        RECT 2.955 1.280 3.340 1.450 ;
        RECT 0.115 0.610 0.445 1.110 ;
        RECT 1.240 0.940 1.630 1.200 ;
        RECT 1.800 1.110 3.340 1.280 ;
        RECT 0.680 0.085 1.010 0.940 ;
        RECT 1.240 0.770 3.005 0.940 ;
        RECT 3.510 0.925 3.680 1.725 ;
        RECT 1.240 0.420 1.630 0.770 ;
        RECT 2.335 0.085 2.665 0.600 ;
        RECT 2.835 0.425 3.005 0.770 ;
        RECT 3.175 0.595 3.680 0.925 ;
        RECT 3.850 1.225 4.150 1.555 ;
        RECT 4.720 1.350 5.020 1.725 ;
        RECT 5.190 1.790 5.440 2.065 ;
        RECT 5.610 1.960 5.940 3.245 ;
        RECT 6.110 1.790 6.440 2.700 ;
        RECT 6.645 1.960 6.975 3.245 ;
        RECT 7.595 2.140 7.925 3.245 ;
        RECT 8.595 2.140 8.925 3.245 ;
        RECT 5.190 1.630 6.935 1.790 ;
        RECT 5.190 1.620 8.595 1.630 ;
        RECT 3.850 0.425 4.020 1.225 ;
        RECT 2.835 0.255 4.020 0.425 ;
        RECT 4.190 0.085 4.440 0.810 ;
        RECT 4.670 0.450 5.000 1.030 ;
        RECT 5.190 0.950 5.360 1.620 ;
        RECT 6.765 1.300 8.595 1.620 ;
        RECT 5.180 0.620 5.360 0.950 ;
        RECT 5.535 0.770 6.725 0.950 ;
        RECT 5.535 0.450 5.785 0.770 ;
        RECT 4.670 0.280 5.785 0.450 ;
        RECT 5.965 0.085 6.295 0.600 ;
        RECT 6.465 0.345 6.725 0.770 ;
        RECT 6.955 0.085 7.215 1.130 ;
        RECT 7.815 0.085 8.145 0.710 ;
        RECT 8.675 0.085 9.005 0.710 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__dlrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.260 0.835 1.930 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.690 1.335 2.150 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.270 1.575 1.280 ;
        RECT 0.005 1.165 2.675 1.270 ;
        RECT 4.690 1.165 8.155 1.240 ;
        RECT 0.005 0.245 8.155 1.165 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
        RECT 4.625 1.580 5.695 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.524500 ;
    PORT
      LAYER li1 ;
        RECT 5.765 1.820 6.130 2.980 ;
        RECT 5.960 1.100 6.130 1.820 ;
        RECT 5.790 0.350 6.130 1.100 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.537600 ;
    PORT
      LAYER li1 ;
        RECT 7.715 0.350 8.050 2.980 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.095 2.100 0.545 2.980 ;
        RECT 0.735 2.320 1.065 3.245 ;
        RECT 1.235 2.560 1.565 2.980 ;
        RECT 2.380 2.730 2.710 3.245 ;
        RECT 1.235 2.390 4.145 2.560 ;
        RECT 1.235 2.320 1.675 2.390 ;
        RECT 0.095 1.090 0.265 2.100 ;
        RECT 1.505 1.520 1.675 2.320 ;
        RECT 1.845 1.880 2.910 2.220 ;
        RECT 3.260 2.050 3.805 2.220 ;
        RECT 2.075 1.710 3.340 1.880 ;
        RECT 1.135 1.260 1.905 1.520 ;
        RECT 0.095 0.750 0.445 1.090 ;
        RECT 1.135 0.920 1.465 1.260 ;
        RECT 2.075 1.090 2.245 1.710 ;
        RECT 1.695 0.920 2.245 1.090 ;
        RECT 2.535 0.750 2.865 1.510 ;
        RECT 0.095 0.580 2.865 0.750 ;
        RECT 3.035 1.470 3.340 1.710 ;
        RECT 3.035 0.505 3.205 1.470 ;
        RECT 3.510 1.300 3.680 2.050 ;
        RECT 3.975 1.800 4.145 2.390 ;
        RECT 4.480 2.060 5.020 3.245 ;
        RECT 5.220 1.890 5.560 2.900 ;
        RECT 6.300 2.100 6.550 3.245 ;
        RECT 3.850 1.470 4.145 1.800 ;
        RECT 4.315 1.720 5.560 1.890 ;
        RECT 4.315 1.470 4.645 1.720 ;
        RECT 5.390 1.600 5.560 1.720 ;
        RECT 6.720 1.630 7.065 2.980 ;
        RECT 7.265 1.820 7.515 3.245 ;
        RECT 4.890 1.300 5.220 1.550 ;
        RECT 3.510 1.130 5.220 1.300 ;
        RECT 5.390 1.270 5.790 1.600 ;
        RECT 6.720 1.300 7.500 1.630 ;
        RECT 3.510 1.055 4.135 1.130 ;
        RECT 3.375 0.725 4.135 1.055 ;
        RECT 5.390 0.960 5.560 1.270 ;
        RECT 0.625 0.085 0.955 0.410 ;
        RECT 2.340 0.085 2.675 0.410 ;
        RECT 3.035 0.255 4.260 0.505 ;
        RECT 4.705 0.085 5.035 0.960 ;
        RECT 5.205 0.350 5.560 0.960 ;
        RECT 6.300 0.085 6.550 1.130 ;
        RECT 6.720 0.540 7.060 1.300 ;
        RECT 7.290 0.085 7.540 1.130 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__dlxbn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.440 1.450 0.815 1.780 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.695 1.315 2.150 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.280 1.575 1.360 ;
        RECT 0.005 1.240 2.135 1.280 ;
        RECT 0.005 1.165 2.610 1.240 ;
        RECT 4.680 1.165 9.115 1.240 ;
        RECT 0.005 0.245 9.115 1.165 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.800 6.590 2.070 ;
        RECT 5.885 1.130 6.115 1.800 ;
        RECT 5.885 0.850 6.505 1.130 ;
        RECT 6.245 0.355 6.505 0.850 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 8.225 1.820 8.555 2.980 ;
        RECT 8.325 1.130 8.495 1.820 ;
        RECT 8.245 0.350 8.495 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.100 2.100 0.445 2.980 ;
        RECT 0.650 2.320 0.980 3.245 ;
        RECT 1.150 2.560 1.485 2.980 ;
        RECT 2.360 2.730 2.690 3.245 ;
        RECT 1.150 2.390 4.275 2.560 ;
        RECT 1.150 2.320 1.655 2.390 ;
        RECT 0.100 1.250 0.270 2.100 ;
        RECT 1.485 1.525 1.655 2.320 ;
        RECT 1.825 1.880 2.155 2.220 ;
        RECT 3.230 2.050 3.935 2.220 ;
        RECT 1.825 1.710 3.385 1.880 ;
        RECT 1.135 1.260 1.885 1.525 ;
        RECT 0.100 0.750 0.445 1.250 ;
        RECT 1.135 0.920 1.465 1.260 ;
        RECT 2.055 1.090 2.225 1.710 ;
        RECT 1.695 0.920 2.225 1.090 ;
        RECT 2.515 0.750 2.845 1.540 ;
        RECT 0.100 0.580 2.845 0.750 ;
        RECT 3.015 1.470 3.385 1.710 ;
        RECT 3.015 0.505 3.185 1.470 ;
        RECT 3.555 1.185 3.725 2.050 ;
        RECT 4.105 1.750 4.275 2.390 ;
        RECT 4.670 2.070 5.080 3.245 ;
        RECT 5.250 2.410 5.655 2.980 ;
        RECT 5.890 2.580 6.140 3.245 ;
        RECT 6.710 2.580 7.040 3.245 ;
        RECT 5.250 2.240 6.955 2.410 ;
        RECT 5.250 1.890 5.655 2.240 ;
        RECT 3.895 1.420 4.275 1.750 ;
        RECT 4.445 1.720 5.655 1.890 ;
        RECT 4.445 1.355 4.775 1.720 ;
        RECT 4.985 1.185 5.315 1.550 ;
        RECT 3.555 1.055 5.315 1.185 ;
        RECT 3.355 1.015 5.315 1.055 ;
        RECT 3.355 0.725 4.070 1.015 ;
        RECT 5.485 0.845 5.655 1.720 ;
        RECT 6.785 1.630 6.955 2.240 ;
        RECT 6.285 1.300 6.955 1.630 ;
        RECT 7.215 1.650 7.545 2.980 ;
        RECT 7.775 1.820 8.025 3.245 ;
        RECT 8.755 1.820 9.005 3.245 ;
        RECT 7.215 1.320 8.155 1.650 ;
        RECT 7.215 1.130 7.515 1.320 ;
        RECT 0.625 0.085 0.955 0.410 ;
        RECT 2.285 0.085 2.640 0.410 ;
        RECT 3.015 0.255 4.265 0.505 ;
        RECT 4.630 0.085 5.015 0.845 ;
        RECT 5.185 0.350 5.655 0.845 ;
        RECT 5.825 0.085 6.075 0.680 ;
        RECT 6.675 0.085 7.005 1.130 ;
        RECT 7.185 0.450 7.515 1.130 ;
        RECT 7.745 0.085 8.075 1.130 ;
        RECT 8.675 0.085 9.005 1.130 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__dlxbn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.220 0.835 1.890 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.180 1.335 1.550 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.735 1.240 2.680 1.280 ;
        RECT 5.690 1.240 7.165 1.260 ;
        RECT 0.010 1.170 2.680 1.240 ;
        RECT 4.410 1.170 8.155 1.240 ;
        RECT 0.010 0.245 8.155 1.170 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.537600 ;
    PORT
      LAYER li1 ;
        RECT 5.765 1.820 6.125 2.980 ;
        RECT 5.955 1.150 6.125 1.820 ;
        RECT 5.795 0.370 6.125 1.150 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.535700 ;
    PORT
      LAYER li1 ;
        RECT 7.715 0.350 8.050 2.980 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.095 2.715 0.440 2.925 ;
        RECT 0.640 2.885 0.970 3.245 ;
        RECT 0.095 2.545 1.760 2.715 ;
        RECT 0.095 2.060 0.440 2.545 ;
        RECT 0.095 1.050 0.265 2.060 ;
        RECT 1.170 1.890 1.420 2.375 ;
        RECT 1.590 2.230 1.760 2.545 ;
        RECT 1.930 2.610 2.180 2.820 ;
        RECT 2.380 2.780 2.710 3.245 ;
        RECT 1.930 2.440 4.100 2.610 ;
        RECT 4.490 2.545 5.035 3.245 ;
        RECT 1.930 2.400 2.180 2.440 ;
        RECT 1.590 2.060 2.875 2.230 ;
        RECT 1.170 1.720 2.330 1.890 ;
        RECT 1.505 1.470 2.330 1.720 ;
        RECT 2.545 1.470 2.875 2.060 ;
        RECT 3.045 1.480 3.215 2.440 ;
        RECT 3.385 1.820 3.555 2.270 ;
        RECT 3.770 2.050 4.100 2.440 ;
        RECT 5.205 2.320 5.535 2.980 ;
        RECT 4.315 1.990 5.535 2.320 ;
        RECT 6.295 2.100 6.545 3.245 ;
        RECT 3.385 1.650 5.035 1.820 ;
        RECT 0.095 0.540 0.450 1.050 ;
        RECT 1.505 1.010 1.675 1.470 ;
        RECT 3.045 1.190 3.515 1.480 ;
        RECT 0.630 0.085 0.960 1.010 ;
        RECT 1.130 0.750 1.675 1.010 ;
        RECT 1.845 1.020 3.515 1.190 ;
        RECT 1.845 0.920 2.175 1.020 ;
        RECT 3.780 0.850 3.950 1.650 ;
        RECT 4.705 1.240 5.035 1.650 ;
        RECT 5.205 1.650 5.535 1.990 ;
        RECT 6.720 1.650 7.050 2.980 ;
        RECT 7.270 1.820 7.520 3.245 ;
        RECT 5.205 1.320 5.775 1.650 ;
        RECT 6.720 1.320 7.320 1.650 ;
        RECT 5.205 1.070 5.375 1.320 ;
        RECT 1.130 0.580 3.080 0.750 ;
        RECT 3.310 0.680 3.950 0.850 ;
        RECT 1.130 0.350 1.675 0.580 ;
        RECT 2.910 0.510 3.080 0.580 ;
        RECT 2.355 0.085 2.740 0.410 ;
        RECT 2.910 0.255 4.075 0.510 ;
        RECT 4.520 0.085 4.850 1.060 ;
        RECT 5.020 0.350 5.375 1.070 ;
        RECT 6.295 0.085 6.545 1.150 ;
        RECT 6.720 0.560 7.055 1.320 ;
        RECT 7.285 0.085 7.535 1.130 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__dlxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.565 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.500 1.315 1.830 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.630 1.255 1.575 1.440 ;
        RECT 0.005 1.240 1.575 1.255 ;
        RECT 3.825 1.240 5.720 1.245 ;
        RECT 0.005 1.165 2.810 1.240 ;
        RECT 3.825 1.165 6.715 1.240 ;
        RECT 0.005 0.245 6.715 1.165 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.545000 ;
    PORT
      LAYER li1 ;
        RECT 6.270 0.350 6.605 2.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.120 1.905 0.450 2.955 ;
        RECT 0.620 2.075 0.950 3.245 ;
        RECT 1.155 2.610 1.655 2.955 ;
        RECT 2.360 2.780 2.705 3.245 ;
        RECT 2.875 2.905 4.180 3.075 ;
        RECT 2.875 2.610 3.045 2.905 ;
        RECT 1.155 2.440 3.045 2.610 ;
        RECT 1.155 2.075 1.655 2.440 ;
        RECT 0.120 1.735 0.775 1.905 ;
        RECT 0.605 1.010 0.775 1.735 ;
        RECT 1.485 1.770 1.655 2.075 ;
        RECT 1.825 1.940 2.225 2.270 ;
        RECT 3.330 2.065 3.840 2.735 ;
        RECT 2.055 1.895 2.225 1.940 ;
        RECT 1.485 1.330 1.885 1.770 ;
        RECT 0.115 0.830 0.775 1.010 ;
        RECT 1.135 1.000 1.885 1.330 ;
        RECT 0.115 0.660 1.315 0.830 ;
        RECT 1.485 0.760 1.885 1.000 ;
        RECT 2.055 1.725 3.500 1.895 ;
        RECT 0.115 0.555 0.445 0.660 ;
        RECT 0.625 0.085 0.955 0.490 ;
        RECT 1.145 0.425 1.315 0.660 ;
        RECT 2.055 0.595 2.305 1.725 ;
        RECT 2.475 1.225 2.970 1.555 ;
        RECT 3.180 1.470 3.500 1.725 ;
        RECT 2.475 0.425 2.645 1.225 ;
        RECT 1.145 0.255 2.645 0.425 ;
        RECT 2.815 0.085 3.145 1.055 ;
        RECT 3.315 0.585 3.485 1.470 ;
        RECT 3.670 1.055 3.840 2.065 ;
        RECT 4.010 1.785 4.180 2.905 ;
        RECT 4.470 2.525 5.065 3.245 ;
        RECT 5.265 2.355 5.655 2.980 ;
        RECT 4.350 2.025 5.655 2.355 ;
        RECT 5.265 1.940 5.655 2.025 ;
        RECT 4.010 1.455 4.340 1.785 ;
        RECT 4.510 1.305 5.315 1.635 ;
        RECT 5.485 1.630 5.655 1.940 ;
        RECT 5.825 1.820 6.075 3.245 ;
        RECT 4.510 1.055 4.680 1.305 ;
        RECT 5.485 1.300 5.885 1.630 ;
        RECT 5.485 1.135 5.655 1.300 ;
        RECT 3.655 0.805 4.680 1.055 ;
        RECT 3.315 0.255 4.355 0.585 ;
        RECT 4.850 0.085 5.100 1.135 ;
        RECT 5.280 0.455 5.655 1.135 ;
        RECT 5.840 0.085 6.090 1.130 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__dlxtn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.450 1.315 1.780 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 1.575 1.280 ;
        RECT 3.845 1.240 5.690 1.245 ;
        RECT 0.005 1.165 2.810 1.240 ;
        RECT 3.845 1.165 7.195 1.240 ;
        RECT 0.005 0.245 7.195 1.165 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
        RECT 4.670 1.635 5.740 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.638000 ;
    PORT
      LAYER li1 ;
        RECT 6.260 1.920 6.635 2.890 ;
        RECT 6.415 1.125 6.585 1.920 ;
        RECT 6.320 0.350 6.585 1.125 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.265 2.120 0.595 2.980 ;
        RECT 0.765 2.290 1.095 3.245 ;
        RECT 1.265 2.610 1.655 2.980 ;
        RECT 2.360 2.780 2.705 3.245 ;
        RECT 2.875 2.905 4.190 3.075 ;
        RECT 2.875 2.610 3.045 2.905 ;
        RECT 1.265 2.440 3.045 2.610 ;
        RECT 0.265 1.950 0.795 2.120 ;
        RECT 1.265 2.100 1.655 2.440 ;
        RECT 0.625 1.130 0.795 1.950 ;
        RECT 1.485 1.770 1.655 2.100 ;
        RECT 1.825 1.970 2.225 2.270 ;
        RECT 3.330 2.140 3.850 2.735 ;
        RECT 1.825 1.940 3.510 1.970 ;
        RECT 2.055 1.800 3.510 1.940 ;
        RECT 1.485 1.170 1.885 1.770 ;
        RECT 0.115 0.750 0.795 1.130 ;
        RECT 1.135 0.920 1.885 1.170 ;
        RECT 1.485 0.760 1.885 0.920 ;
        RECT 0.115 0.580 1.315 0.750 ;
        RECT 2.055 0.595 2.305 1.800 ;
        RECT 2.475 1.300 2.970 1.630 ;
        RECT 3.180 1.470 3.510 1.800 ;
        RECT 1.145 0.425 1.315 0.580 ;
        RECT 2.475 0.425 2.645 1.300 ;
        RECT 0.625 0.085 0.955 0.410 ;
        RECT 1.145 0.255 2.645 0.425 ;
        RECT 2.815 0.085 3.145 1.055 ;
        RECT 3.315 0.585 3.485 1.470 ;
        RECT 3.680 1.055 3.850 2.140 ;
        RECT 4.020 1.815 4.190 2.905 ;
        RECT 4.360 2.625 5.080 3.245 ;
        RECT 5.250 2.355 5.580 2.955 ;
        RECT 4.360 2.025 5.580 2.355 ;
        RECT 5.250 1.965 5.580 2.025 ;
        RECT 4.020 1.485 4.350 1.815 ;
        RECT 5.250 1.795 5.675 1.965 ;
        RECT 5.845 1.820 6.060 3.245 ;
        RECT 6.835 1.820 7.085 3.245 ;
        RECT 5.505 1.625 5.675 1.795 ;
        RECT 4.990 1.315 5.335 1.625 ;
        RECT 4.080 1.295 5.335 1.315 ;
        RECT 5.505 1.295 6.245 1.625 ;
        RECT 4.080 1.145 5.160 1.295 ;
        RECT 4.080 1.055 4.250 1.145 ;
        RECT 5.505 1.125 5.675 1.295 ;
        RECT 3.655 0.805 4.250 1.055 ;
        RECT 3.315 0.255 4.375 0.585 ;
        RECT 4.820 0.085 5.150 0.975 ;
        RECT 5.330 0.955 5.675 1.125 ;
        RECT 5.330 0.355 5.580 0.955 ;
        RECT 5.845 0.085 6.140 1.125 ;
        RECT 6.755 0.085 7.085 1.130 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__dlxtn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.500 1.315 1.830 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.630 1.255 1.575 1.440 ;
        RECT 0.005 1.240 1.575 1.255 ;
        RECT 0.005 1.165 2.810 1.240 ;
        RECT 5.760 1.165 8.155 1.240 ;
        RECT 0.005 0.245 8.155 1.165 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.270300 ;
    PORT
      LAYER li1 ;
        RECT 6.315 1.990 6.645 2.980 ;
        RECT 7.315 2.150 7.545 2.980 ;
        RECT 7.315 1.990 8.035 2.150 ;
        RECT 6.315 1.820 8.035 1.990 ;
        RECT 7.805 1.150 8.035 1.820 ;
        RECT 6.265 0.980 8.035 1.150 ;
        RECT 6.265 0.350 6.615 0.980 ;
        RECT 7.295 0.350 7.545 0.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.135 2.120 0.465 2.980 ;
        RECT 0.635 2.290 0.965 3.245 ;
        RECT 1.135 2.560 1.655 2.980 ;
        RECT 2.360 2.730 2.820 3.245 ;
        RECT 2.990 2.905 4.220 3.075 ;
        RECT 2.990 2.560 3.160 2.905 ;
        RECT 1.135 2.390 3.160 2.560 ;
        RECT 0.135 1.950 0.795 2.120 ;
        RECT 1.135 2.100 1.655 2.390 ;
        RECT 0.625 1.130 0.795 1.950 ;
        RECT 1.485 1.770 1.655 2.100 ;
        RECT 1.825 1.940 2.225 2.220 ;
        RECT 3.360 2.060 3.880 2.735 ;
        RECT 2.055 1.890 2.225 1.940 ;
        RECT 1.485 1.330 1.885 1.770 ;
        RECT 0.115 0.830 0.795 1.130 ;
        RECT 1.135 1.000 1.885 1.330 ;
        RECT 0.115 0.660 1.315 0.830 ;
        RECT 1.485 0.760 1.885 1.000 ;
        RECT 2.055 1.720 3.540 1.890 ;
        RECT 0.115 0.555 0.445 0.660 ;
        RECT 0.625 0.085 0.955 0.490 ;
        RECT 1.145 0.425 1.315 0.660 ;
        RECT 2.055 0.595 2.305 1.720 ;
        RECT 2.475 1.220 3.000 1.550 ;
        RECT 3.210 1.470 3.540 1.720 ;
        RECT 2.475 0.425 2.645 1.220 ;
        RECT 1.145 0.255 2.645 0.425 ;
        RECT 2.815 0.085 3.145 1.050 ;
        RECT 3.315 0.505 3.485 1.470 ;
        RECT 3.710 1.055 3.880 2.060 ;
        RECT 4.050 1.735 4.220 2.905 ;
        RECT 4.390 2.590 5.145 3.245 ;
        RECT 5.315 2.305 5.645 2.980 ;
        RECT 4.390 1.990 5.645 2.305 ;
        RECT 5.815 2.160 6.145 3.245 ;
        RECT 6.815 2.160 7.145 3.245 ;
        RECT 7.715 2.320 8.045 3.245 ;
        RECT 4.390 1.975 5.830 1.990 ;
        RECT 5.315 1.820 5.830 1.975 ;
        RECT 4.050 1.405 4.380 1.735 ;
        RECT 5.660 1.650 5.830 1.820 ;
        RECT 4.550 1.320 5.490 1.650 ;
        RECT 5.660 1.320 7.490 1.650 ;
        RECT 4.550 1.055 4.720 1.320 ;
        RECT 5.660 1.150 5.830 1.320 ;
        RECT 3.655 0.725 4.720 1.055 ;
        RECT 3.315 0.255 4.445 0.505 ;
        RECT 4.890 0.085 5.140 1.055 ;
        RECT 5.320 0.980 5.830 1.150 ;
        RECT 5.320 0.375 5.570 0.980 ;
        RECT 5.750 0.085 6.080 0.810 ;
        RECT 6.785 0.085 7.115 0.810 ;
        RECT 7.715 0.085 8.045 0.810 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__dlxtn_4

#--------EOF---------

MACRO sky130_fd_sc_hs__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.595 1.850 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.350 6.715 1.780 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.145 1.280 4.005 1.295 ;
        RECT 1.145 1.120 7.675 1.280 ;
        RECT 0.005 0.245 7.675 1.120 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
        RECT 4.110 1.505 5.865 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 7.230 1.820 7.595 2.980 ;
        RECT 7.425 1.150 7.595 1.820 ;
        RECT 7.235 0.390 7.595 1.150 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.115 2.100 0.445 3.245 ;
        RECT 0.645 2.100 0.945 2.980 ;
        RECT 0.775 1.770 0.945 2.100 ;
        RECT 1.125 2.785 1.455 2.980 ;
        RECT 1.660 2.955 1.995 3.245 ;
        RECT 2.165 2.785 2.970 2.985 ;
        RECT 1.125 2.735 2.970 2.785 ;
        RECT 3.140 2.845 4.040 3.015 ;
        RECT 4.840 2.845 5.170 3.245 ;
        RECT 1.125 2.615 2.335 2.735 ;
        RECT 1.125 1.940 1.455 2.615 ;
        RECT 3.140 2.565 3.310 2.845 ;
        RECT 5.340 2.675 6.525 2.700 ;
        RECT 2.505 2.445 3.310 2.565 ;
        RECT 2.080 2.395 3.310 2.445 ;
        RECT 3.590 2.505 6.525 2.675 ;
        RECT 2.080 2.275 2.675 2.395 ;
        RECT 2.080 1.940 2.330 2.275 ;
        RECT 2.845 2.105 3.420 2.225 ;
        RECT 2.515 2.055 3.420 2.105 ;
        RECT 2.515 1.935 3.015 2.055 ;
        RECT 0.775 1.100 1.165 1.770 ;
        RECT 1.335 1.355 2.345 1.525 ;
        RECT 0.775 1.010 0.945 1.100 ;
        RECT 0.115 0.085 0.445 1.010 ;
        RECT 0.615 0.420 0.945 1.010 ;
        RECT 1.335 0.930 1.505 1.355 ;
        RECT 1.175 0.405 1.505 0.930 ;
        RECT 1.675 0.085 2.005 1.185 ;
        RECT 2.175 0.925 2.345 1.355 ;
        RECT 2.515 1.265 2.685 1.935 ;
        RECT 3.590 1.885 3.760 2.505 ;
        RECT 3.185 1.765 3.760 1.885 ;
        RECT 2.855 1.715 3.760 1.765 ;
        RECT 3.930 2.165 5.625 2.335 ;
        RECT 2.855 1.435 3.355 1.715 ;
        RECT 3.930 1.545 4.100 2.165 ;
        RECT 4.270 1.665 4.815 1.995 ;
        RECT 3.525 1.275 4.100 1.545 ;
        RECT 2.515 1.105 3.355 1.265 ;
        RECT 2.515 1.095 4.395 1.105 ;
        RECT 3.015 0.935 4.395 1.095 ;
        RECT 2.175 0.765 2.845 0.925 ;
        RECT 4.065 0.775 4.395 0.935 ;
        RECT 2.175 0.755 3.895 0.765 ;
        RECT 2.675 0.595 3.895 0.755 ;
        RECT 4.565 0.750 4.815 1.665 ;
        RECT 5.375 1.170 5.625 2.165 ;
        RECT 5.845 1.950 6.525 2.505 ;
        RECT 6.730 1.950 7.060 3.245 ;
        RECT 5.845 1.350 6.175 1.950 ;
        RECT 6.005 1.170 6.175 1.350 ;
        RECT 6.895 1.320 7.255 1.650 ;
        RECT 5.375 0.920 5.835 1.170 ;
        RECT 6.005 0.920 6.410 1.170 ;
        RECT 6.895 0.750 7.065 1.320 ;
        RECT 2.175 0.425 2.505 0.585 ;
        RECT 4.565 0.580 7.065 0.750 ;
        RECT 4.565 0.425 4.815 0.580 ;
        RECT 2.175 0.255 4.815 0.425 ;
        RECT 4.995 0.085 5.325 0.410 ;
        RECT 6.590 0.085 7.055 0.410 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__dlxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlygate4sd1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.895 0.920 3.675 1.240 ;
        RECT 0.010 0.245 3.675 0.920 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.509700 ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.815 3.740 3.060 ;
        RECT 3.450 1.120 3.740 1.815 ;
        RECT 3.325 0.355 3.740 1.120 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.395 1.720 2.725 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.610 1.720 2.395 ;
        RECT 1.985 1.995 2.345 2.190 ;
        RECT 2.825 2.165 3.155 3.245 ;
        RECT 1.985 1.825 3.155 1.995 ;
        RECT 2.910 1.625 3.155 1.825 ;
        RECT 1.475 1.380 2.740 1.610 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.635 1.720 1.380 ;
        RECT 2.910 1.295 3.280 1.625 ;
        RECT 2.910 1.210 3.155 1.295 ;
        RECT 1.985 1.040 3.155 1.210 ;
        RECT 1.985 0.710 2.345 1.040 ;
        RECT 1.415 0.305 1.720 0.635 ;
        RECT 2.825 0.085 3.155 0.870 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__dlygate4sd1_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlygate4sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlygate4sd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.895 0.920 3.675 1.240 ;
        RECT 0.010 0.245 3.675 0.920 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.509700 ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.815 3.740 3.060 ;
        RECT 3.450 1.120 3.740 1.815 ;
        RECT 3.325 0.355 3.740 1.120 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.395 1.720 2.725 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.610 1.720 2.395 ;
        RECT 1.985 1.995 2.345 2.190 ;
        RECT 2.825 2.165 3.155 3.245 ;
        RECT 1.985 1.825 3.155 1.995 ;
        RECT 2.910 1.625 3.155 1.825 ;
        RECT 1.475 1.380 2.740 1.610 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.635 1.720 1.380 ;
        RECT 2.910 1.295 3.280 1.625 ;
        RECT 2.910 1.210 3.155 1.295 ;
        RECT 1.985 1.040 3.155 1.210 ;
        RECT 1.985 0.710 2.345 1.040 ;
        RECT 1.415 0.305 1.720 0.635 ;
        RECT 2.825 0.085 3.155 0.870 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__dlygate4sd2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlygate4sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlygate4sd3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.190 0.730 1.860 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.895 0.920 3.675 1.240 ;
        RECT 0.010 0.245 3.675 0.920 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.509700 ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.815 3.740 3.060 ;
        RECT 3.450 1.120 3.740 1.815 ;
        RECT 3.325 0.355 3.740 1.120 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.095 2.205 0.400 2.725 ;
        RECT 0.575 2.380 0.905 3.245 ;
        RECT 1.415 2.395 1.720 2.725 ;
        RECT 0.095 2.030 1.305 2.205 ;
        RECT 0.975 1.020 1.305 2.030 ;
        RECT 0.095 0.820 1.305 1.020 ;
        RECT 1.475 1.610 1.720 2.395 ;
        RECT 1.985 1.995 2.345 2.190 ;
        RECT 2.825 2.165 3.155 3.245 ;
        RECT 1.985 1.825 3.155 1.995 ;
        RECT 2.910 1.625 3.155 1.825 ;
        RECT 1.475 1.380 2.740 1.610 ;
        RECT 0.095 0.305 0.410 0.820 ;
        RECT 0.585 0.085 0.915 0.650 ;
        RECT 1.475 0.635 1.720 1.380 ;
        RECT 2.910 1.295 3.280 1.625 ;
        RECT 2.910 1.210 3.155 1.295 ;
        RECT 1.985 1.040 3.155 1.210 ;
        RECT 1.985 0.710 2.345 1.040 ;
        RECT 1.415 0.305 1.720 0.635 ;
        RECT 2.825 0.085 3.155 0.870 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__dlygate4sd3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlymetal6s2s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlymetal6s2s_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.355 0.555 1.765 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 4.320 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER met1 ;
        RECT 0.965 2.320 4.210 2.490 ;
        RECT 0.965 1.920 1.345 2.320 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.590 2.310 0.885 3.245 ;
        RECT 0.100 2.140 0.430 2.225 ;
        RECT 0.100 1.935 0.895 2.140 ;
        RECT 0.725 1.605 0.895 1.935 ;
        RECT 1.065 1.835 1.380 3.075 ;
        RECT 2.100 2.310 2.395 3.245 ;
        RECT 1.550 2.140 1.870 2.225 ;
        RECT 2.565 2.160 2.865 3.075 ;
        RECT 3.585 2.310 3.880 3.245 ;
        RECT 1.550 1.895 2.335 2.140 ;
        RECT 1.210 1.605 1.380 1.835 ;
        RECT 2.165 1.605 2.335 1.895 ;
        RECT 2.505 1.835 2.865 2.160 ;
        RECT 3.070 2.140 3.400 2.225 ;
        RECT 4.050 2.160 4.350 3.075 ;
        RECT 3.070 1.895 3.805 2.140 ;
        RECT 2.695 1.605 2.865 1.835 ;
        RECT 3.605 1.605 3.805 1.895 ;
        RECT 3.975 1.835 4.350 2.160 ;
        RECT 0.725 1.275 1.040 1.605 ;
        RECT 1.210 1.315 1.995 1.605 ;
        RECT 0.725 1.145 0.895 1.275 ;
        RECT 0.100 0.975 0.895 1.145 ;
        RECT 1.210 1.075 1.380 1.315 ;
        RECT 2.165 1.275 2.525 1.605 ;
        RECT 2.695 1.315 3.435 1.605 ;
        RECT 2.165 1.145 2.335 1.275 ;
        RECT 0.100 0.700 0.395 0.975 ;
        RECT 0.590 0.085 0.920 0.805 ;
        RECT 1.090 0.255 1.380 1.075 ;
        RECT 1.550 0.975 2.335 1.145 ;
        RECT 2.695 1.075 2.865 1.315 ;
        RECT 3.605 1.275 4.010 1.605 ;
        RECT 3.605 1.145 3.775 1.275 ;
        RECT 1.550 0.700 1.835 0.975 ;
        RECT 2.030 0.085 2.360 0.805 ;
        RECT 2.530 0.255 2.865 1.075 ;
        RECT 3.060 0.975 3.775 1.145 ;
        RECT 4.180 1.075 4.350 1.835 ;
        RECT 3.060 0.700 3.275 0.975 ;
        RECT 3.470 0.085 3.800 0.805 ;
        RECT 3.970 0.255 4.350 1.075 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 2.555 1.950 2.725 2.120 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
      LAYER met1 ;
        RECT 2.405 1.920 2.785 2.150 ;
        RECT 3.845 1.920 4.225 2.150 ;
  END
END sky130_fd_sc_hs__dlymetal6s2s_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlymetal6s4s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlymetal6s4s_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.355 0.555 1.765 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 4.320 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER met1 ;
        RECT 0.965 2.320 4.210 2.490 ;
        RECT 2.405 1.920 2.785 2.320 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.590 2.310 0.885 3.245 ;
        RECT 0.100 2.140 0.430 2.225 ;
        RECT 0.100 1.935 0.895 2.140 ;
        RECT 0.725 1.605 0.895 1.935 ;
        RECT 1.065 1.835 1.380 3.075 ;
        RECT 2.100 2.310 2.395 3.245 ;
        RECT 1.550 2.140 1.870 2.225 ;
        RECT 2.565 2.160 2.865 3.075 ;
        RECT 3.585 2.310 3.880 3.245 ;
        RECT 1.550 1.895 2.335 2.140 ;
        RECT 1.210 1.605 1.380 1.835 ;
        RECT 2.165 1.605 2.335 1.895 ;
        RECT 2.505 1.835 2.865 2.160 ;
        RECT 3.070 2.140 3.400 2.225 ;
        RECT 4.050 2.160 4.350 3.075 ;
        RECT 3.070 1.895 3.805 2.140 ;
        RECT 2.695 1.605 2.865 1.835 ;
        RECT 3.605 1.605 3.805 1.895 ;
        RECT 3.975 1.835 4.350 2.160 ;
        RECT 0.725 1.275 1.040 1.605 ;
        RECT 1.210 1.315 1.995 1.605 ;
        RECT 0.725 1.145 0.895 1.275 ;
        RECT 0.100 0.975 0.895 1.145 ;
        RECT 1.210 1.075 1.380 1.315 ;
        RECT 2.165 1.275 2.525 1.605 ;
        RECT 2.695 1.315 3.435 1.605 ;
        RECT 2.165 1.145 2.335 1.275 ;
        RECT 0.100 0.700 0.395 0.975 ;
        RECT 0.590 0.085 0.920 0.805 ;
        RECT 1.090 0.255 1.380 1.075 ;
        RECT 1.550 0.975 2.335 1.145 ;
        RECT 2.695 1.075 2.865 1.315 ;
        RECT 3.605 1.275 4.010 1.605 ;
        RECT 3.605 1.145 3.775 1.275 ;
        RECT 1.550 0.700 1.835 0.975 ;
        RECT 2.030 0.085 2.360 0.805 ;
        RECT 2.530 0.255 2.865 1.075 ;
        RECT 3.060 0.975 3.775 1.145 ;
        RECT 4.180 1.075 4.350 1.835 ;
        RECT 3.060 0.700 3.275 0.975 ;
        RECT 3.470 0.085 3.800 0.805 ;
        RECT 3.970 0.255 4.350 1.075 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 2.555 1.950 2.725 2.120 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
      LAYER met1 ;
        RECT 0.965 1.920 1.345 2.150 ;
        RECT 3.845 1.920 4.225 2.150 ;
  END
END sky130_fd_sc_hs__dlymetal6s4s_1

#--------EOF---------

MACRO sky130_fd_sc_hs__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dlymetal6s6s_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.355 0.555 1.765 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.245 4.320 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER met1 ;
        RECT 0.965 2.320 4.225 2.490 ;
        RECT 3.845 1.920 4.225 2.320 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.590 2.310 0.885 3.245 ;
        RECT 0.100 2.140 0.430 2.225 ;
        RECT 0.100 1.935 0.895 2.140 ;
        RECT 0.725 1.605 0.895 1.935 ;
        RECT 1.065 1.835 1.380 3.075 ;
        RECT 2.100 2.310 2.395 3.245 ;
        RECT 1.550 2.140 1.870 2.225 ;
        RECT 2.565 2.160 2.865 3.075 ;
        RECT 3.585 2.310 3.880 3.245 ;
        RECT 1.550 1.895 2.335 2.140 ;
        RECT 1.210 1.605 1.380 1.835 ;
        RECT 2.165 1.605 2.335 1.895 ;
        RECT 2.505 1.835 2.865 2.160 ;
        RECT 3.070 2.140 3.400 2.225 ;
        RECT 4.050 2.160 4.350 3.075 ;
        RECT 3.070 1.895 3.805 2.140 ;
        RECT 2.695 1.605 2.865 1.835 ;
        RECT 3.605 1.605 3.805 1.895 ;
        RECT 3.975 1.835 4.350 2.160 ;
        RECT 0.725 1.275 1.040 1.605 ;
        RECT 1.210 1.315 1.995 1.605 ;
        RECT 0.725 1.145 0.895 1.275 ;
        RECT 0.100 0.975 0.895 1.145 ;
        RECT 1.210 1.075 1.380 1.315 ;
        RECT 2.165 1.275 2.525 1.605 ;
        RECT 2.695 1.315 3.435 1.605 ;
        RECT 2.165 1.145 2.335 1.275 ;
        RECT 0.100 0.700 0.395 0.975 ;
        RECT 0.590 0.085 0.920 0.805 ;
        RECT 1.090 0.255 1.380 1.075 ;
        RECT 1.550 0.975 2.335 1.145 ;
        RECT 2.695 1.075 2.865 1.315 ;
        RECT 3.605 1.275 4.010 1.605 ;
        RECT 3.605 1.145 3.775 1.275 ;
        RECT 1.550 0.700 1.835 0.975 ;
        RECT 2.030 0.085 2.360 0.805 ;
        RECT 2.530 0.255 2.865 1.075 ;
        RECT 3.060 0.975 3.775 1.145 ;
        RECT 4.180 1.075 4.350 1.835 ;
        RECT 3.060 0.700 3.275 0.975 ;
        RECT 3.470 0.085 3.800 0.805 ;
        RECT 3.970 0.255 4.350 1.075 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 1.115 1.950 1.285 2.120 ;
        RECT 2.555 1.950 2.725 2.120 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
      LAYER met1 ;
        RECT 0.965 1.920 1.345 2.150 ;
        RECT 2.405 1.920 2.785 2.150 ;
  END
END sky130_fd_sc_hs__dlymetal6s6s_1

#--------EOF---------

MACRO sky130_fd_sc_hs__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ebufn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.500 1.795 1.830 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.376500 ;
    PORT
      LAYER li1 ;
        RECT 1.865 2.590 2.195 3.010 ;
        RECT 0.665 2.420 2.195 2.590 ;
        RECT 0.665 1.830 0.835 2.420 ;
        RECT 1.865 2.340 2.195 2.420 ;
        RECT 0.425 1.500 0.835 1.830 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.280 1.050 3.650 1.240 ;
        RECT 0.130 0.245 3.650 1.050 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.235 1.820 3.755 2.980 ;
        RECT 3.585 1.130 3.755 1.820 ;
        RECT 3.210 0.350 3.755 1.130 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.085 2.000 0.445 2.880 ;
        RECT 0.650 2.760 0.980 3.245 ;
        RECT 1.185 2.170 1.695 2.250 ;
        RECT 1.185 2.000 2.135 2.170 ;
        RECT 2.365 2.050 2.695 3.245 ;
        RECT 0.085 1.320 0.255 2.000 ;
        RECT 1.965 1.880 2.135 2.000 ;
        RECT 1.965 1.710 3.065 1.880 ;
        RECT 2.460 1.650 3.065 1.710 ;
        RECT 1.870 1.320 2.200 1.340 ;
        RECT 0.085 1.150 2.200 1.320 ;
        RECT 2.460 1.320 3.415 1.650 ;
        RECT 0.085 0.455 0.530 1.150 ;
        RECT 2.460 0.980 2.660 1.320 ;
        RECT 0.700 0.085 0.985 0.850 ;
        RECT 1.155 0.810 2.660 0.980 ;
        RECT 1.155 0.455 1.450 0.810 ;
        RECT 2.390 0.085 2.720 0.640 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__ebufn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ebufn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 3.865 1.780 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.582000 ;
    PORT
      LAYER li1 ;
        RECT 2.965 1.180 3.295 1.650 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 2.415 1.240 ;
        RECT 0.005 0.245 4.280 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.599200 ;
    PORT
      LAYER li1 ;
        RECT 0.645 2.150 0.975 2.735 ;
        RECT 0.645 1.970 1.795 2.150 ;
        RECT 0.535 1.800 1.795 1.970 ;
        RECT 0.535 1.130 0.705 1.800 ;
        RECT 0.535 0.615 0.875 1.130 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.145 2.905 1.475 3.075 ;
        RECT 1.680 2.920 2.010 3.245 ;
        RECT 0.145 2.140 0.475 2.905 ;
        RECT 1.145 2.750 1.475 2.905 ;
        RECT 2.215 2.750 2.545 2.980 ;
        RECT 1.145 2.580 2.545 2.750 ;
        RECT 3.225 2.610 3.705 3.245 ;
        RECT 1.145 2.320 1.475 2.580 ;
        RECT 3.875 2.410 4.205 2.860 ;
        RECT 1.965 2.240 4.205 2.410 ;
        RECT 1.965 1.630 2.135 2.240 ;
        RECT 0.875 1.300 2.135 1.630 ;
        RECT 2.395 1.820 3.105 2.070 ;
        RECT 3.875 1.950 4.205 2.240 ;
        RECT 0.115 0.425 0.365 1.130 ;
        RECT 1.045 0.960 2.225 1.130 ;
        RECT 1.045 0.425 1.375 0.960 ;
        RECT 0.115 0.255 1.375 0.425 ;
        RECT 1.545 0.085 1.795 0.790 ;
        RECT 1.975 0.350 2.225 0.960 ;
        RECT 2.395 1.010 2.725 1.820 ;
        RECT 4.035 1.030 4.205 1.950 ;
        RECT 2.395 0.325 3.170 1.010 ;
        RECT 3.340 0.085 3.670 1.010 ;
        RECT 3.840 0.350 4.205 1.030 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__ebufn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ebufn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.300 0.805 1.780 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.951000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.180 1.285 1.550 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.101200 ;
    PORT
      LAYER li1 ;
        RECT 3.970 1.990 4.300 2.735 ;
        RECT 4.870 1.990 5.205 2.735 ;
        RECT 3.970 1.820 5.205 1.990 ;
        RECT 5.035 1.150 5.205 1.820 ;
        RECT 4.015 0.980 5.205 1.150 ;
        RECT 4.015 0.595 4.345 0.980 ;
        RECT 4.875 0.595 5.205 0.980 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.085 2.560 0.365 2.980 ;
        RECT 0.565 2.730 0.920 3.245 ;
        RECT 1.800 2.570 1.970 2.820 ;
        RECT 2.170 2.740 2.500 3.245 ;
        RECT 2.700 2.570 2.870 2.980 ;
        RECT 0.085 2.390 1.630 2.560 ;
        RECT 1.800 2.400 2.870 2.570 ;
        RECT 0.085 1.950 0.365 2.390 ;
        RECT 1.460 2.230 1.630 2.390 ;
        RECT 0.085 1.130 0.255 1.950 ;
        RECT 1.040 1.890 1.290 2.220 ;
        RECT 1.460 2.060 2.530 2.230 ;
        RECT 1.040 1.720 1.775 1.890 ;
        RECT 0.085 0.350 0.405 1.130 ;
        RECT 1.455 1.010 1.775 1.720 ;
        RECT 2.360 1.650 2.530 2.060 ;
        RECT 2.700 1.990 2.870 2.400 ;
        RECT 3.070 2.160 3.320 3.245 ;
        RECT 3.520 2.905 5.650 3.075 ;
        RECT 3.520 1.990 3.770 2.905 ;
        RECT 4.470 2.160 4.700 2.905 ;
        RECT 2.700 1.820 3.770 1.990 ;
        RECT 5.400 1.820 5.650 2.905 ;
        RECT 2.360 1.480 4.830 1.650 ;
        RECT 3.820 1.320 4.830 1.480 ;
        RECT 0.585 0.085 0.915 1.010 ;
        RECT 1.095 0.300 1.775 1.010 ;
        RECT 1.945 1.150 2.975 1.310 ;
        RECT 1.945 1.140 3.835 1.150 ;
        RECT 1.945 0.350 2.115 1.140 ;
        RECT 2.805 0.980 3.835 1.140 ;
        RECT 2.295 0.085 2.625 0.970 ;
        RECT 2.805 0.350 2.975 0.980 ;
        RECT 3.155 0.085 3.405 0.810 ;
        RECT 3.585 0.425 3.835 0.980 ;
        RECT 4.525 0.425 4.695 0.810 ;
        RECT 5.405 0.425 5.655 1.130 ;
        RECT 3.585 0.255 5.655 0.425 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__ebufn_4

#--------EOF---------

MACRO sky130_fd_sc_hs__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ebufn_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 9.645 1.180 9.975 1.550 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.623000 ;
    PORT
      LAYER li1 ;
        RECT 8.265 1.180 9.475 1.550 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.560 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 7.740 1.240 ;
        RECT 8.710 0.245 10.555 1.240 ;
        RECT 0.000 0.000 10.560 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.750 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.560 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.360500 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.990 0.900 2.735 ;
        RECT 1.520 1.990 1.850 2.735 ;
        RECT 2.420 1.990 2.750 2.735 ;
        RECT 3.370 1.990 3.700 2.735 ;
        RECT 0.545 1.820 3.700 1.990 ;
        RECT 0.545 1.150 0.835 1.820 ;
        RECT 0.545 0.980 3.760 1.150 ;
        RECT 0.545 0.595 0.875 0.980 ;
        RECT 1.430 0.595 1.760 0.980 ;
        RECT 2.430 0.595 2.760 0.980 ;
        RECT 3.430 0.595 3.760 0.980 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.560 3.415 ;
        RECT 0.120 2.905 4.200 3.075 ;
        RECT 0.120 1.820 0.370 2.905 ;
        RECT 1.085 2.160 1.350 2.905 ;
        RECT 2.050 2.160 2.220 2.905 ;
        RECT 2.920 2.160 3.190 2.905 ;
        RECT 3.870 2.560 4.200 2.905 ;
        RECT 4.370 2.730 4.700 3.245 ;
        RECT 4.870 2.560 5.200 2.980 ;
        RECT 5.370 2.730 5.700 3.245 ;
        RECT 5.870 2.560 6.200 2.980 ;
        RECT 6.370 2.730 6.700 3.245 ;
        RECT 6.870 2.730 7.200 2.980 ;
        RECT 7.405 2.900 7.735 3.245 ;
        RECT 7.940 2.730 8.270 2.980 ;
        RECT 6.870 2.560 8.270 2.730 ;
        RECT 9.165 2.560 9.495 3.245 ;
        RECT 3.870 2.390 7.200 2.560 ;
        RECT 9.665 2.390 9.945 2.980 ;
        RECT 7.585 2.220 9.945 2.390 ;
        RECT 3.870 2.050 7.755 2.220 ;
        RECT 3.870 1.650 4.040 2.050 ;
        RECT 1.035 1.480 4.040 1.650 ;
        RECT 7.925 1.800 9.045 2.050 ;
        RECT 9.665 1.890 9.945 2.220 ;
        RECT 10.115 2.060 10.445 3.245 ;
        RECT 1.035 1.320 3.655 1.480 ;
        RECT 4.720 1.310 7.550 1.470 ;
        RECT 3.940 1.300 7.550 1.310 ;
        RECT 3.940 1.140 5.050 1.300 ;
        RECT 0.115 0.425 0.365 1.130 ;
        RECT 1.055 0.425 1.225 0.810 ;
        RECT 1.930 0.425 2.260 0.810 ;
        RECT 2.930 0.425 3.260 0.810 ;
        RECT 3.940 0.425 4.110 1.140 ;
        RECT 0.115 0.255 4.110 0.425 ;
        RECT 4.290 0.085 4.620 0.970 ;
        RECT 4.800 0.350 5.050 1.140 ;
        RECT 5.230 0.085 5.400 1.130 ;
        RECT 5.580 0.350 5.830 1.300 ;
        RECT 6.010 0.085 6.260 1.130 ;
        RECT 6.440 0.350 6.690 1.300 ;
        RECT 6.870 0.085 7.120 1.130 ;
        RECT 7.300 0.350 7.550 1.300 ;
        RECT 7.925 1.010 8.095 1.800 ;
        RECT 9.665 1.720 10.315 1.890 ;
        RECT 10.145 1.010 10.315 1.720 ;
        RECT 7.925 0.670 9.150 1.010 ;
        RECT 7.720 0.340 9.150 0.670 ;
        RECT 9.330 0.085 9.500 1.010 ;
        RECT 9.680 0.840 10.315 1.010 ;
        RECT 9.680 0.340 9.930 0.840 ;
        RECT 10.110 0.085 10.445 0.600 ;
        RECT 0.000 -0.085 10.560 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
  END
END sky130_fd_sc_hs__ebufn_8

#--------EOF---------

MACRO sky130_fd_sc_hs__edfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__edfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.715 1.180 4.385 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.980 0.835 1.990 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.285000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.450 1.905 1.780 ;
    END
  END DE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.525 1.035 5.435 1.240 ;
        RECT 8.470 1.140 9.775 1.240 ;
        RECT 12.655 1.140 14.395 1.260 ;
        RECT 7.395 1.035 14.395 1.140 ;
        RECT 3.525 0.920 14.395 1.035 ;
        RECT 0.005 0.245 14.395 0.920 ;
        RECT 0.000 0.000 14.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.590 3.520 ;
        RECT 4.945 1.650 6.045 1.660 ;
        RECT 11.870 1.645 12.940 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.400 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 12.925 1.820 13.340 2.980 ;
        RECT 12.925 1.000 13.095 1.820 ;
        RECT 12.765 0.620 13.095 1.000 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 13.990 1.820 14.315 2.980 ;
        RECT 14.145 1.150 14.315 1.820 ;
        RECT 13.955 0.370 14.315 1.150 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.400 3.415 ;
        RECT 0.085 2.460 0.445 2.980 ;
        RECT 0.955 2.630 1.205 3.245 ;
        RECT 1.375 2.905 2.225 3.075 ;
        RECT 1.375 2.460 1.545 2.905 ;
        RECT 0.085 2.290 1.545 2.460 ;
        RECT 0.085 0.750 0.255 2.290 ;
        RECT 1.715 2.120 1.885 2.735 ;
        RECT 2.055 2.460 2.225 2.905 ;
        RECT 2.395 2.630 2.645 3.245 ;
        RECT 3.155 2.480 3.545 2.960 ;
        RECT 3.715 2.650 4.045 3.245 ;
        RECT 5.105 2.650 5.435 3.245 ;
        RECT 5.605 2.890 6.445 3.060 ;
        RECT 5.605 2.480 5.775 2.890 ;
        RECT 6.650 2.720 6.980 2.980 ;
        RECT 7.695 2.885 8.025 3.245 ;
        RECT 3.155 2.460 5.775 2.480 ;
        RECT 2.055 2.310 5.775 2.460 ;
        RECT 6.550 2.550 6.980 2.720 ;
        RECT 8.195 2.755 9.405 2.925 ;
        RECT 8.195 2.715 8.365 2.755 ;
        RECT 2.055 2.290 3.545 2.310 ;
        RECT 1.005 1.950 2.665 2.120 ;
        RECT 1.005 1.280 1.335 1.950 ;
        RECT 1.005 1.110 2.000 1.280 ;
        RECT 0.085 0.420 0.600 0.750 ;
        RECT 1.090 0.085 1.420 0.810 ;
        RECT 1.650 0.480 2.000 1.110 ;
        RECT 2.335 0.980 2.665 1.950 ;
        RECT 2.875 0.980 3.205 1.990 ;
        RECT 3.375 0.810 3.545 2.290 ;
        RECT 4.165 1.810 4.965 2.140 ;
        RECT 4.555 1.010 4.725 1.810 ;
        RECT 5.215 1.470 5.385 2.310 ;
        RECT 5.955 2.140 6.355 2.380 ;
        RECT 5.555 1.970 6.355 2.140 ;
        RECT 5.555 1.810 6.125 1.970 ;
        RECT 5.215 1.300 5.785 1.470 ;
        RECT 2.170 0.085 2.500 0.810 ;
        RECT 3.000 0.350 3.545 0.810 ;
        RECT 3.715 0.085 3.885 1.010 ;
        RECT 4.065 0.840 4.725 1.010 ;
        RECT 4.065 0.350 4.395 0.840 ;
        RECT 4.585 0.085 4.915 0.670 ;
        RECT 5.095 0.425 5.345 1.130 ;
        RECT 5.535 0.595 5.785 1.300 ;
        RECT 5.955 0.425 6.125 1.810 ;
        RECT 6.550 1.910 6.720 2.550 ;
        RECT 7.150 2.545 8.365 2.715 ;
        RECT 7.150 2.380 7.320 2.545 ;
        RECT 6.890 2.080 7.320 2.380 ;
        RECT 8.700 2.375 9.030 2.585 ;
        RECT 8.230 2.125 9.030 2.375 ;
        RECT 7.930 1.910 8.260 1.955 ;
        RECT 6.550 1.740 8.260 1.910 ;
        RECT 6.550 1.685 6.720 1.740 ;
        RECT 6.295 1.515 6.720 1.685 ;
        RECT 7.930 1.645 8.260 1.740 ;
        RECT 6.295 0.595 6.465 1.515 ;
        RECT 7.205 1.475 7.535 1.570 ;
        RECT 8.700 1.475 9.030 2.125 ;
        RECT 9.235 1.790 9.405 2.755 ;
        RECT 9.575 1.960 9.905 3.245 ;
        RECT 10.445 2.155 10.775 2.980 ;
        RECT 11.495 2.325 12.280 3.245 ;
        RECT 10.445 1.985 11.445 2.155 ;
        RECT 12.450 2.120 12.700 2.845 ;
        RECT 9.235 1.620 10.625 1.790 ;
        RECT 6.635 1.135 6.885 1.345 ;
        RECT 7.205 1.305 9.030 1.475 ;
        RECT 10.295 1.460 10.625 1.620 ;
        RECT 6.635 0.965 7.810 1.135 ;
        RECT 6.635 0.425 6.885 0.965 ;
        RECT 5.095 0.255 6.885 0.425 ;
        RECT 7.220 0.085 7.470 0.795 ;
        RECT 7.640 0.425 7.810 0.965 ;
        RECT 7.980 0.595 8.150 1.305 ;
        RECT 9.200 1.290 10.085 1.450 ;
        RECT 10.835 1.290 11.105 1.800 ;
        RECT 9.200 1.135 11.105 1.290 ;
        RECT 8.320 1.120 11.105 1.135 ;
        RECT 11.275 1.485 11.445 1.985 ;
        RECT 11.615 1.805 12.700 2.120 ;
        RECT 13.540 1.820 13.790 3.245 ;
        RECT 11.615 1.725 12.485 1.805 ;
        RECT 11.275 1.155 11.985 1.485 ;
        RECT 8.320 0.965 9.370 1.120 ;
        RECT 8.320 0.425 8.490 0.965 ;
        RECT 11.275 0.950 11.445 1.155 ;
        RECT 7.640 0.255 8.490 0.425 ;
        RECT 8.660 0.085 8.910 0.770 ;
        RECT 9.540 0.620 11.445 0.950 ;
        RECT 11.655 0.085 11.985 0.985 ;
        RECT 12.155 0.425 12.485 1.725 ;
        RECT 13.265 1.320 13.975 1.650 ;
        RECT 13.265 0.425 13.435 1.320 ;
        RECT 12.155 0.255 13.435 0.425 ;
        RECT 13.605 0.085 13.775 1.150 ;
        RECT 0.000 -0.085 14.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 3.035 1.580 3.205 1.750 ;
        RECT 12.155 1.580 12.325 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
      LAYER met1 ;
        RECT 2.975 1.735 3.265 1.780 ;
        RECT 12.095 1.735 12.385 1.780 ;
        RECT 2.975 1.595 12.385 1.735 ;
        RECT 2.975 1.550 3.265 1.595 ;
        RECT 12.095 1.550 12.385 1.595 ;
  END
END sky130_fd_sc_hs__edfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__edfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__edfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.450 1.180 3.780 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.980 0.805 1.990 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.285000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.110 1.845 1.440 ;
    END
  END DE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.250 1.000 5.205 1.240 ;
        RECT 8.420 1.220 9.890 1.240 ;
        RECT 7.345 1.000 9.890 1.220 ;
        RECT 3.250 0.985 9.890 1.000 ;
        RECT 1.465 0.920 9.890 0.985 ;
        RECT 11.905 0.920 12.955 1.240 ;
        RECT 0.090 0.245 12.955 0.920 ;
        RECT 0.000 0.000 12.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.150 3.520 ;
        RECT 3.525 1.580 4.590 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.960 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518900 ;
    PORT
      LAYER li1 ;
        RECT 12.075 1.550 12.405 2.980 ;
        RECT 12.075 1.130 12.345 1.550 ;
        RECT 12.015 0.350 12.345 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.085 2.350 0.435 2.980 ;
        RECT 0.945 2.520 1.195 3.245 ;
        RECT 1.365 2.905 2.215 3.075 ;
        RECT 1.365 2.350 1.535 2.905 ;
        RECT 0.085 2.180 1.535 2.350 ;
        RECT 0.085 0.810 0.255 2.180 ;
        RECT 0.975 1.780 1.305 2.010 ;
        RECT 1.705 1.780 1.875 2.735 ;
        RECT 2.045 2.120 2.215 2.905 ;
        RECT 2.385 2.290 2.635 3.245 ;
        RECT 3.670 2.650 4.000 3.245 ;
        RECT 5.020 2.650 5.270 3.245 ;
        RECT 5.995 2.690 6.245 2.980 ;
        RECT 3.100 2.480 3.475 2.620 ;
        RECT 5.440 2.520 6.245 2.690 ;
        RECT 6.415 2.520 6.775 2.980 ;
        RECT 7.410 2.750 7.740 3.245 ;
        RECT 8.505 2.750 8.835 3.245 ;
        RECT 5.440 2.480 5.610 2.520 ;
        RECT 3.100 2.310 5.610 2.480 ;
        RECT 3.100 2.120 3.475 2.310 ;
        RECT 2.045 1.950 3.270 2.120 ;
        RECT 0.975 1.610 2.385 1.780 ;
        RECT 0.975 0.940 1.305 1.610 ;
        RECT 2.055 1.385 2.385 1.610 ;
        RECT 2.555 1.045 2.930 1.780 ;
        RECT 0.085 0.340 0.530 0.810 ;
        RECT 0.975 0.770 1.820 0.940 ;
        RECT 3.100 0.875 3.270 1.950 ;
        RECT 3.950 1.470 4.900 2.140 ;
        RECT 5.130 1.650 5.300 2.310 ;
        RECT 5.825 2.140 6.245 2.300 ;
        RECT 5.470 1.970 6.245 2.140 ;
        RECT 5.470 1.820 5.995 1.970 ;
        RECT 5.130 1.480 5.655 1.650 ;
        RECT 3.950 1.010 4.120 1.470 ;
        RECT 1.020 0.085 1.350 0.600 ;
        RECT 1.570 0.415 1.820 0.770 ;
        RECT 2.000 0.085 2.330 0.875 ;
        RECT 2.790 0.415 3.270 0.875 ;
        RECT 3.440 0.085 3.610 1.010 ;
        RECT 3.790 0.350 4.120 1.010 ;
        RECT 4.335 0.085 4.585 1.130 ;
        RECT 4.765 0.425 5.095 1.130 ;
        RECT 5.325 0.595 5.655 1.480 ;
        RECT 5.825 0.425 5.995 1.820 ;
        RECT 6.415 1.800 6.585 2.520 ;
        RECT 6.945 2.410 9.800 2.580 ;
        RECT 6.945 2.330 7.115 2.410 ;
        RECT 6.755 2.000 7.115 2.330 ;
        RECT 7.945 2.070 8.440 2.240 ;
        RECT 7.700 1.800 8.030 1.830 ;
        RECT 6.165 1.630 8.030 1.800 ;
        RECT 6.165 0.765 6.335 1.630 ;
        RECT 7.700 1.615 8.030 1.630 ;
        RECT 8.270 1.605 8.440 2.070 ;
        RECT 9.630 1.725 9.800 2.410 ;
        RECT 9.970 2.095 10.220 3.000 ;
        RECT 10.845 2.525 11.385 3.245 ;
        RECT 11.555 2.320 11.885 2.950 ;
        RECT 10.665 2.095 11.885 2.320 ;
        RECT 9.970 1.925 10.405 2.095 ;
        RECT 10.235 1.755 10.945 1.925 ;
        RECT 7.130 1.445 7.460 1.460 ;
        RECT 8.270 1.445 8.940 1.605 ;
        RECT 6.505 1.105 6.960 1.310 ;
        RECT 7.130 1.275 8.940 1.445 ;
        RECT 9.110 1.375 9.460 1.550 ;
        RECT 9.630 1.545 10.065 1.725 ;
        RECT 10.275 1.375 10.605 1.585 ;
        RECT 6.505 0.935 7.760 1.105 ;
        RECT 6.165 0.595 6.620 0.765 ;
        RECT 6.790 0.425 6.960 0.935 ;
        RECT 4.765 0.255 6.960 0.425 ;
        RECT 7.170 0.085 7.420 0.765 ;
        RECT 7.590 0.425 7.760 0.935 ;
        RECT 7.930 0.595 8.100 1.275 ;
        RECT 9.110 1.205 10.605 1.375 ;
        RECT 10.775 1.335 10.945 1.755 ;
        RECT 11.645 1.550 11.885 2.095 ;
        RECT 12.605 1.820 12.855 3.245 ;
        RECT 9.110 1.105 9.280 1.205 ;
        RECT 8.270 0.935 9.280 1.105 ;
        RECT 10.775 1.005 11.505 1.335 ;
        RECT 8.270 0.425 8.440 0.935 ;
        RECT 9.450 0.835 10.945 1.005 ;
        RECT 7.590 0.255 8.440 0.425 ;
        RECT 8.610 0.085 8.860 0.765 ;
        RECT 9.450 0.350 9.780 0.835 ;
        RECT 11.675 0.810 11.845 1.550 ;
        RECT 10.350 0.085 11.310 0.665 ;
        RECT 11.490 0.335 11.845 0.810 ;
        RECT 12.515 0.085 12.845 1.130 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 2.555 1.580 2.725 1.750 ;
        RECT 11.675 1.580 11.845 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
      LAYER met1 ;
        RECT 2.495 1.735 2.785 1.780 ;
        RECT 11.615 1.735 11.905 1.780 ;
        RECT 2.495 1.595 11.905 1.735 ;
        RECT 2.495 1.550 2.785 1.595 ;
        RECT 11.615 1.550 11.905 1.595 ;
  END
END sky130_fd_sc_hs__edfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 1.975 1.780 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.327000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.760 1.315 1.780 ;
        RECT 0.455 1.430 1.315 1.760 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.325 1.370 1.275 1.450 ;
        RECT 0.325 0.245 2.210 1.370 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.950 2.315 2.980 ;
        RECT 2.145 1.180 2.315 1.950 ;
        RECT 1.770 0.480 2.315 1.180 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.390 2.100 0.720 2.580 ;
        RECT 0.110 1.930 0.720 2.100 ;
        RECT 0.925 1.950 1.255 3.245 ;
        RECT 0.110 1.250 0.280 1.930 ;
        RECT 0.110 0.560 0.770 1.250 ;
        RECT 0.110 0.255 0.780 0.560 ;
        RECT 0.950 0.085 1.280 1.260 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__einvn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 0.810 3.255 1.550 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.120 0.550 2.130 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.025 0.920 3.265 1.240 ;
        RECT 0.020 0.790 3.265 0.920 ;
        RECT 0.020 0.245 3.315 0.790 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.546900 ;
    PORT
      LAYER li1 ;
        RECT 2.465 1.820 2.795 2.735 ;
        RECT 2.465 1.130 2.755 1.820 ;
        RECT 2.425 0.770 2.755 1.130 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.110 2.300 0.360 3.245 ;
        RECT 0.560 2.300 0.890 2.980 ;
        RECT 0.720 1.650 0.890 2.300 ;
        RECT 1.115 1.990 1.400 2.980 ;
        RECT 1.580 2.160 1.815 3.245 ;
        RECT 2.015 2.905 3.245 3.075 ;
        RECT 2.015 1.990 2.295 2.905 ;
        RECT 1.115 1.820 2.295 1.990 ;
        RECT 2.965 1.820 3.245 2.905 ;
        RECT 0.720 1.320 1.160 1.650 ;
        RECT 0.720 0.810 0.890 1.320 ;
        RECT 0.130 0.085 0.380 0.810 ;
        RECT 0.560 0.350 0.890 0.810 ;
        RECT 1.135 0.980 2.245 1.150 ;
        RECT 1.135 0.350 1.385 0.980 ;
        RECT 1.565 0.085 1.895 0.790 ;
        RECT 2.075 0.600 2.245 0.980 ;
        RECT 2.075 0.350 3.200 0.600 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__einvn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__einvn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.035 1.180 5.155 1.550 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.951000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.275 1.240 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.890 3.815 2.735 ;
        RECT 4.385 1.890 4.715 2.735 ;
        RECT 3.485 1.720 4.715 1.890 ;
        RECT 3.485 1.550 3.815 1.720 ;
        RECT 3.615 1.130 3.815 1.550 ;
        RECT 3.615 1.010 3.865 1.130 ;
        RECT 3.615 0.770 4.655 1.010 ;
        RECT 4.485 0.595 4.655 0.770 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.175 1.950 0.425 3.245 ;
        RECT 0.625 1.310 0.955 2.980 ;
        RECT 1.185 1.650 1.435 2.980 ;
        RECT 1.635 1.820 1.885 3.245 ;
        RECT 2.085 1.650 2.335 2.980 ;
        RECT 2.535 1.820 2.865 3.245 ;
        RECT 3.035 2.905 5.165 3.075 ;
        RECT 3.035 1.650 3.285 2.905 ;
        RECT 4.015 2.060 4.185 2.905 ;
        RECT 4.915 1.820 5.165 2.905 ;
        RECT 1.185 1.480 3.285 1.650 ;
        RECT 0.625 1.130 1.295 1.310 ;
        RECT 0.115 0.085 0.365 1.130 ;
        RECT 0.545 0.300 1.295 1.130 ;
        RECT 1.465 1.140 3.435 1.310 ;
        RECT 1.465 0.350 1.635 1.140 ;
        RECT 1.815 0.085 2.145 0.970 ;
        RECT 2.325 0.350 2.495 1.140 ;
        RECT 2.675 0.085 3.005 0.970 ;
        RECT 3.185 0.600 3.435 1.140 ;
        RECT 3.185 0.425 4.305 0.600 ;
        RECT 4.835 0.425 5.165 1.010 ;
        RECT 3.185 0.255 5.165 0.425 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__einvn_4

#--------EOF---------

MACRO sky130_fd_sc_hs__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvn_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.232000 ;
    PORT
      LAYER li1 ;
        RECT 5.995 1.350 8.995 1.780 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.623000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.630 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.065 0.245 9.115 1.240 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.332400 ;
    PORT
      LAYER li1 ;
        RECT 5.555 2.120 5.725 2.735 ;
        RECT 6.425 2.120 6.755 2.735 ;
        RECT 7.325 2.120 7.655 2.735 ;
        RECT 8.225 2.120 8.555 2.735 ;
        RECT 5.555 1.950 8.555 2.120 ;
        RECT 5.555 1.780 5.725 1.950 ;
        RECT 4.925 1.550 5.725 1.780 ;
        RECT 5.455 1.130 5.725 1.550 ;
        RECT 6.315 1.130 8.505 1.180 ;
        RECT 5.455 1.010 8.505 1.130 ;
        RECT 5.455 0.770 6.645 1.010 ;
        RECT 7.325 0.615 7.495 1.010 ;
        RECT 8.175 0.615 8.505 1.010 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.115 1.820 0.445 3.245 ;
        RECT 0.615 1.335 0.945 2.980 ;
        RECT 1.175 1.835 1.425 2.980 ;
        RECT 1.625 2.005 1.955 3.245 ;
        RECT 2.125 1.835 2.375 2.980 ;
        RECT 2.575 2.005 2.905 3.245 ;
        RECT 3.075 1.835 3.325 2.980 ;
        RECT 3.525 2.005 3.855 3.245 ;
        RECT 4.025 2.120 4.355 2.980 ;
        RECT 4.525 2.290 4.855 3.245 ;
        RECT 5.025 2.905 9.005 3.075 ;
        RECT 5.025 2.120 5.355 2.905 ;
        RECT 5.925 2.290 6.255 2.905 ;
        RECT 6.955 2.290 7.125 2.905 ;
        RECT 7.855 2.290 8.025 2.905 ;
        RECT 4.025 1.950 5.355 2.120 ;
        RECT 8.755 1.950 9.005 2.905 ;
        RECT 4.025 1.835 4.495 1.950 ;
        RECT 1.175 1.665 4.495 1.835 ;
        RECT 1.525 1.380 4.415 1.470 ;
        RECT 0.615 1.130 1.355 1.335 ;
        RECT 0.175 0.085 0.505 0.990 ;
        RECT 0.685 0.325 1.355 1.130 ;
        RECT 1.525 1.300 5.275 1.380 ;
        RECT 1.525 0.350 1.695 1.300 ;
        RECT 1.875 0.085 2.125 1.130 ;
        RECT 2.305 0.350 2.555 1.300 ;
        RECT 2.735 0.085 3.065 1.130 ;
        RECT 3.235 0.350 3.485 1.300 ;
        RECT 4.165 1.210 5.275 1.300 ;
        RECT 3.665 0.085 3.995 1.130 ;
        RECT 4.165 0.350 4.415 1.210 ;
        RECT 4.595 0.085 4.925 1.040 ;
        RECT 5.105 0.600 5.275 1.210 ;
        RECT 6.815 0.600 7.145 0.825 ;
        RECT 5.105 0.425 7.145 0.600 ;
        RECT 7.675 0.425 8.005 0.825 ;
        RECT 8.675 0.425 9.005 1.130 ;
        RECT 5.105 0.255 9.005 0.425 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__einvn_8

#--------EOF---------

MACRO sky130_fd_sc_hs__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.300 2.275 1.780 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.440 1.315 1.780 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.045 0.920 2.395 1.240 ;
        RECT 0.200 0.245 2.395 0.920 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.505900 ;
    PORT
      LAYER li1 ;
        RECT 1.955 2.275 2.285 2.980 ;
        RECT 1.605 1.950 2.285 2.275 ;
        RECT 1.605 1.130 1.775 1.950 ;
        RECT 1.605 0.960 2.285 1.130 ;
        RECT 1.955 0.350 2.285 0.960 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.105 2.745 0.890 3.075 ;
        RECT 0.105 2.010 0.880 2.745 ;
        RECT 1.085 2.020 1.415 3.245 ;
        RECT 0.105 1.060 0.275 2.010 ;
        RECT 0.105 0.410 0.940 1.060 ;
        RECT 1.135 0.085 1.420 1.130 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__einvp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__einvp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 2.480 0.260 2.810 0.670 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.360 1.240 3.355 1.250 ;
        RECT 0.050 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.180 0.920 2.735 ;
        RECT 0.670 0.625 0.920 1.180 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.905 1.265 3.075 ;
        RECT 0.115 1.820 0.365 2.905 ;
        RECT 1.095 1.650 1.265 2.905 ;
        RECT 1.465 1.820 1.715 3.245 ;
        RECT 1.915 1.650 2.165 2.980 ;
        RECT 1.095 1.480 2.165 1.650 ;
        RECT 1.100 1.140 2.210 1.310 ;
        RECT 0.160 0.425 0.490 1.010 ;
        RECT 1.100 0.425 1.270 1.140 ;
        RECT 0.160 0.255 1.270 0.425 ;
        RECT 1.450 0.085 1.780 0.970 ;
        RECT 1.950 0.350 2.210 1.140 ;
        RECT 2.415 1.140 2.745 2.980 ;
        RECT 2.915 2.300 3.245 3.245 ;
        RECT 2.415 0.840 2.800 1.140 ;
        RECT 2.980 0.085 3.245 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__einvp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.430 1.780 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.723000 ;
    PORT
      LAYER li1 ;
        RECT 4.980 1.300 5.650 1.630 ;
        RECT 5.405 1.180 5.650 1.300 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.615 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.221900 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 0.945 2.735 ;
        RECT 1.565 2.120 1.895 2.735 ;
        RECT 0.615 1.950 1.895 2.120 ;
        RECT 1.615 1.180 1.895 1.950 ;
        RECT 0.615 1.010 1.945 1.180 ;
        RECT 0.615 0.660 0.945 1.010 ;
        RECT 1.615 0.660 1.945 1.010 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 2.905 2.395 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 1.115 2.290 1.365 2.905 ;
        RECT 2.065 1.810 2.395 2.905 ;
        RECT 2.565 1.980 2.815 3.245 ;
        RECT 3.015 1.810 3.265 2.980 ;
        RECT 3.465 1.980 3.725 3.245 ;
        RECT 4.395 2.980 4.785 2.990 ;
        RECT 3.925 1.810 4.175 2.980 ;
        RECT 2.065 1.640 4.175 1.810 ;
        RECT 4.395 1.820 5.195 2.980 ;
        RECT 5.395 1.820 5.645 3.245 ;
        RECT 4.395 1.640 4.785 1.820 ;
        RECT 2.115 1.300 4.445 1.470 ;
        RECT 0.115 0.425 0.445 1.130 ;
        RECT 1.115 0.425 1.445 0.800 ;
        RECT 2.115 0.425 2.445 1.300 ;
        RECT 0.115 0.255 2.445 0.425 ;
        RECT 2.615 0.085 2.945 1.130 ;
        RECT 3.115 0.350 3.445 1.300 ;
        RECT 3.615 0.085 3.945 1.130 ;
        RECT 4.115 0.350 4.445 1.300 ;
        RECT 4.615 1.130 4.785 1.640 ;
        RECT 4.615 0.350 5.005 1.130 ;
        RECT 5.175 0.085 5.505 1.010 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__einvp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__einvp_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.232000 ;
    PORT
      LAYER li1 ;
        RECT 0.410 1.180 3.460 1.550 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.167000 ;
    PORT
      LAYER li1 ;
        RECT 8.435 1.410 8.765 1.550 ;
        RECT 8.435 1.180 8.995 1.410 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 9.045 1.240 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.328200 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.890 0.890 2.735 ;
        RECT 1.460 1.890 1.790 2.735 ;
        RECT 2.360 1.890 2.690 2.735 ;
        RECT 3.260 1.890 3.590 2.735 ;
        RECT 0.560 1.720 4.195 1.890 ;
        RECT 3.705 1.550 4.195 1.720 ;
        RECT 3.705 1.010 3.875 1.550 ;
        RECT 0.625 0.840 3.875 1.010 ;
        RECT 0.625 0.615 0.875 0.840 ;
        RECT 1.545 0.615 1.875 0.840 ;
        RECT 2.545 0.615 2.875 0.840 ;
        RECT 3.545 0.595 3.875 0.840 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.110 2.905 3.960 3.075 ;
        RECT 0.110 1.820 0.375 2.905 ;
        RECT 1.070 2.060 1.275 2.905 ;
        RECT 1.970 2.060 2.190 2.905 ;
        RECT 2.875 2.060 3.075 2.905 ;
        RECT 3.790 2.230 3.960 2.905 ;
        RECT 4.160 2.400 4.490 3.245 ;
        RECT 4.690 2.230 4.940 2.980 ;
        RECT 3.790 2.060 4.940 2.230 ;
        RECT 4.690 1.720 4.940 2.060 ;
        RECT 5.140 1.890 5.310 3.245 ;
        RECT 5.510 1.720 5.760 2.980 ;
        RECT 5.960 1.890 6.210 3.245 ;
        RECT 6.410 1.720 6.660 2.980 ;
        RECT 6.860 1.890 7.110 3.245 ;
        RECT 7.310 1.720 7.560 2.980 ;
        RECT 8.235 2.965 8.565 2.980 ;
        RECT 4.690 1.550 7.560 1.720 ;
        RECT 7.775 1.820 8.565 2.965 ;
        RECT 8.765 1.820 9.015 3.245 ;
        RECT 7.775 1.615 8.225 1.820 ;
        RECT 4.055 1.210 7.885 1.380 ;
        RECT 0.115 0.425 0.445 1.010 ;
        RECT 1.045 0.425 1.375 0.670 ;
        RECT 2.045 0.425 2.375 0.670 ;
        RECT 3.045 0.425 3.375 0.670 ;
        RECT 4.055 0.425 4.225 1.210 ;
        RECT 0.115 0.255 4.225 0.425 ;
        RECT 4.405 0.085 4.735 1.040 ;
        RECT 4.905 0.350 5.155 1.210 ;
        RECT 5.335 0.085 5.665 1.040 ;
        RECT 5.845 0.350 6.015 1.210 ;
        RECT 6.195 0.085 6.525 1.040 ;
        RECT 6.705 0.350 6.955 1.210 ;
        RECT 7.125 0.085 7.455 1.040 ;
        RECT 7.635 0.350 7.885 1.210 ;
        RECT 8.055 1.010 8.225 1.615 ;
        RECT 8.055 0.350 8.505 1.010 ;
        RECT 8.675 0.085 8.935 1.010 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__einvp_8

#--------EOF---------

MACRO sky130_fd_sc_hs__fa_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fa_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 0.885 1.220 1.215 1.540 ;
        RECT 1.045 1.090 1.215 1.220 ;
        RECT 3.300 1.090 3.630 1.455 ;
        RECT 4.380 1.105 4.710 1.455 ;
        RECT 5.810 1.320 6.210 1.575 ;
        RECT 5.810 1.105 5.980 1.320 ;
        RECT 4.380 1.090 5.980 1.105 ;
        RECT 1.045 0.935 5.980 1.090 ;
        RECT 1.045 0.920 4.710 0.935 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 6.800 1.320 7.470 1.780 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.738000 ;
    PORT
      LAYER met1 ;
        RECT 1.535 1.735 1.825 1.780 ;
        RECT 3.935 1.735 4.225 1.780 ;
        RECT 4.895 1.735 5.185 1.780 ;
        RECT 1.535 1.595 5.185 1.735 ;
        RECT 1.535 1.550 1.825 1.595 ;
        RECT 3.935 1.550 4.225 1.595 ;
        RECT 4.895 1.550 5.185 1.595 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.145 0.950 1.240 ;
        RECT 7.690 1.145 8.635 1.240 ;
        RECT 0.005 0.245 8.635 1.145 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
        RECT 1.500 1.555 7.480 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.519000 ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.130 8.540 2.980 ;
        RECT 8.210 0.350 8.540 1.130 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.355 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.365 1.130 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.555 2.050 0.885 3.245 ;
        RECT 2.080 2.120 2.410 2.755 ;
        RECT 1.055 1.950 2.410 2.120 ;
        RECT 2.610 2.460 2.860 2.755 ;
        RECT 3.080 2.630 3.410 3.245 ;
        RECT 3.600 2.460 3.930 2.755 ;
        RECT 2.610 2.290 3.930 2.460 ;
        RECT 4.105 2.305 4.435 3.245 ;
        RECT 2.610 1.965 2.860 2.290 ;
        RECT 5.070 2.120 5.495 2.755 ;
        RECT 1.055 1.880 1.225 1.950 ;
        RECT 0.535 1.710 1.225 1.880 ;
        RECT 0.535 1.630 0.705 1.710 ;
        RECT 0.425 1.300 0.705 1.630 ;
        RECT 0.535 0.750 0.705 1.300 ;
        RECT 1.565 1.575 1.795 1.780 ;
        RECT 2.080 1.745 2.410 1.950 ;
        RECT 3.030 1.950 5.495 2.120 ;
        RECT 5.665 2.255 5.950 2.755 ;
        RECT 6.120 2.500 6.825 3.245 ;
        RECT 7.000 2.255 7.320 2.830 ;
        RECT 5.665 2.085 7.320 2.255 ;
        RECT 6.990 1.950 7.320 2.085 ;
        RECT 3.030 1.795 3.200 1.950 ;
        RECT 2.580 1.625 3.200 1.795 ;
        RECT 5.325 1.915 5.495 1.950 ;
        RECT 2.580 1.575 2.750 1.625 ;
        RECT 1.565 1.260 2.115 1.575 ;
        RECT 2.325 1.260 2.750 1.575 ;
        RECT 3.840 1.260 4.195 1.780 ;
        RECT 4.925 1.575 5.155 1.780 ;
        RECT 5.325 1.745 6.550 1.915 ;
        RECT 7.755 1.820 8.085 3.245 ;
        RECT 4.925 1.275 5.640 1.575 ;
        RECT 6.380 1.150 6.550 1.745 ;
        RECT 7.710 1.150 8.040 1.550 ;
        RECT 6.150 0.980 8.040 1.150 ;
        RECT 6.150 0.765 6.320 0.980 ;
        RECT 0.535 0.580 2.270 0.750 ;
        RECT 0.625 0.085 0.980 0.410 ;
        RECT 1.940 0.355 2.270 0.580 ;
        RECT 2.480 0.580 3.910 0.750 ;
        RECT 2.480 0.420 2.890 0.580 ;
        RECT 3.580 0.420 3.910 0.580 ;
        RECT 3.070 0.085 3.400 0.410 ;
        RECT 4.080 0.085 4.555 0.710 ;
        RECT 5.045 0.595 6.320 0.765 ;
        RECT 6.490 0.640 7.590 0.810 ;
        RECT 5.045 0.435 5.375 0.595 ;
        RECT 6.490 0.425 6.660 0.640 ;
        RECT 7.260 0.480 7.590 0.640 ;
        RECT 5.555 0.255 6.660 0.425 ;
        RECT 6.830 0.085 7.080 0.470 ;
        RECT 7.780 0.085 8.030 0.770 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 1.595 1.580 1.765 1.750 ;
        RECT 3.995 1.580 4.165 1.750 ;
        RECT 4.955 1.580 5.125 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__fa_1

#--------EOF---------

MACRO sky130_fd_sc_hs__fa_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fa_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.044000 ;
    PORT
      LAYER met1 ;
        RECT 0.095 1.735 0.385 1.780 ;
        RECT 2.495 1.735 2.785 1.780 ;
        RECT 3.935 1.735 4.225 1.780 ;
        RECT 6.335 1.735 6.625 1.780 ;
        RECT 0.095 1.595 6.625 1.735 ;
        RECT 0.095 1.550 0.385 1.595 ;
        RECT 2.495 1.550 2.785 1.595 ;
        RECT 3.935 1.550 4.225 1.595 ;
        RECT 6.335 1.550 6.625 1.595 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.044000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.920 0.835 2.150 ;
        RECT 0.665 1.575 0.835 1.920 ;
        RECT 0.665 1.245 1.165 1.575 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.783000 ;
    PORT
      LAYER li1 ;
        RECT 3.375 2.120 4.195 2.150 ;
        RECT 2.055 2.105 4.195 2.120 ;
        RECT 2.055 1.950 4.535 2.105 ;
        RECT 2.055 1.575 2.225 1.950 ;
        RECT 3.375 1.935 4.535 1.950 ;
        RECT 3.375 1.575 3.545 1.935 ;
        RECT 4.365 1.915 4.535 1.935 ;
        RECT 4.365 1.745 5.635 1.915 ;
        RECT 1.715 1.260 2.225 1.575 ;
        RECT 3.215 1.260 3.545 1.575 ;
        RECT 5.305 1.260 5.635 1.745 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 9.115 1.265 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
        RECT 0.635 1.555 5.915 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.649600 ;
    PORT
      LAYER li1 ;
        RECT 6.985 1.820 7.555 2.150 ;
        RECT 7.385 1.085 7.555 1.820 ;
        RECT 7.105 0.915 7.555 1.085 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 8.220 1.820 8.575 2.980 ;
        RECT 8.405 1.150 8.575 1.820 ;
        RECT 8.245 0.375 8.575 1.150 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.095 2.490 0.445 2.910 ;
        RECT 0.615 2.660 1.010 3.245 ;
        RECT 1.215 2.490 1.545 2.755 ;
        RECT 0.095 2.320 1.545 2.490 ;
        RECT 0.095 1.950 0.425 2.320 ;
        RECT 1.215 2.085 1.545 2.320 ;
        RECT 1.715 2.290 2.185 2.620 ;
        RECT 2.825 2.290 3.155 3.245 ;
        RECT 3.405 2.490 3.735 2.755 ;
        RECT 3.905 2.660 4.290 3.245 ;
        RECT 4.495 2.490 4.825 2.755 ;
        RECT 3.405 2.320 4.825 2.490 ;
        RECT 1.715 1.915 1.885 2.290 ;
        RECT 4.495 2.275 4.825 2.320 ;
        RECT 5.005 2.490 5.335 2.755 ;
        RECT 6.535 2.660 6.865 3.245 ;
        RECT 7.530 2.730 8.050 3.245 ;
        RECT 5.005 2.320 8.050 2.490 ;
        RECT 5.005 2.085 5.335 2.320 ;
        RECT 0.105 1.300 0.435 1.780 ;
        RECT 1.375 1.745 1.885 1.915 ;
        RECT 0.115 1.075 0.445 1.130 ;
        RECT 1.375 1.090 1.545 1.745 ;
        RECT 2.525 1.575 2.755 1.780 ;
        RECT 3.965 1.575 4.195 1.765 ;
        RECT 2.525 1.260 3.005 1.575 ;
        RECT 3.965 1.260 4.525 1.575 ;
        RECT 4.765 1.090 5.095 1.575 ;
        RECT 6.265 1.350 6.595 1.780 ;
        RECT 7.880 1.650 8.050 2.320 ;
        RECT 8.750 1.820 9.000 3.245 ;
        RECT 6.765 1.255 7.165 1.585 ;
        RECT 7.880 1.320 8.235 1.650 ;
        RECT 6.765 1.090 6.935 1.255 ;
        RECT 0.115 0.905 1.205 1.075 ;
        RECT 1.375 0.920 6.935 1.090 ;
        RECT 0.115 0.375 0.445 0.905 ;
        RECT 1.035 0.750 1.205 0.905 ;
        RECT 0.615 0.085 0.865 0.735 ;
        RECT 1.035 0.420 1.810 0.750 ;
        RECT 1.980 0.375 2.310 0.920 ;
        RECT 2.800 0.085 3.310 0.705 ;
        RECT 3.480 0.580 4.970 0.750 ;
        RECT 3.480 0.375 3.810 0.580 ;
        RECT 4.500 0.420 4.970 0.580 ;
        RECT 5.140 0.745 5.470 0.750 ;
        RECT 7.880 0.745 8.050 1.320 ;
        RECT 5.140 0.575 8.050 0.745 ;
        RECT 3.990 0.085 4.320 0.410 ;
        RECT 5.140 0.375 5.470 0.575 ;
        RECT 6.470 0.085 6.925 0.405 ;
        RECT 7.615 0.085 8.065 0.405 ;
        RECT 8.755 0.085 9.005 1.155 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 1.580 0.325 1.750 ;
        RECT 2.555 1.580 2.725 1.750 ;
        RECT 3.995 1.580 4.165 1.750 ;
        RECT 6.395 1.580 6.565 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__fa_2

#--------EOF---------

MACRO sky130_fd_sc_hs__fa_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fa_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.044000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.245 0.835 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.044000 ;
    PORT
      LAYER li1 ;
        RECT 1.665 1.950 2.650 2.120 ;
        RECT 1.665 1.575 1.835 1.950 ;
        RECT 1.345 1.260 1.835 1.575 ;
        RECT 2.480 1.915 2.650 1.950 ;
        RECT 2.480 1.890 4.620 1.915 ;
        RECT 2.480 1.780 6.085 1.890 ;
        RECT 2.480 1.745 6.595 1.780 ;
        RECT 2.480 1.245 2.810 1.745 ;
        RECT 3.950 1.260 4.280 1.745 ;
        RECT 4.450 1.720 6.595 1.745 ;
        RECT 5.915 1.550 6.595 1.720 ;
        RECT 5.915 1.260 6.340 1.550 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.783000 ;
    PORT
      LAYER met1 ;
        RECT 2.015 1.365 2.305 1.410 ;
        RECT 2.975 1.365 3.265 1.410 ;
        RECT 5.375 1.365 5.665 1.410 ;
        RECT 2.015 1.225 5.665 1.365 ;
        RECT 2.015 1.180 2.305 1.225 ;
        RECT 2.975 1.180 3.265 1.225 ;
        RECT 5.375 1.180 5.665 1.225 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.760 1.240 11.035 1.280 ;
        RECT 0.005 0.245 11.035 1.240 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
        RECT 0.635 1.555 6.620 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 9.145 1.990 9.475 2.980 ;
        RECT 10.095 1.990 10.435 2.980 ;
        RECT 9.145 1.820 10.435 1.990 ;
        RECT 10.165 1.550 10.435 1.820 ;
        RECT 10.165 1.150 10.425 1.550 ;
        RECT 9.305 0.980 10.425 1.150 ;
        RECT 9.305 0.390 9.555 0.980 ;
        RECT 10.165 0.390 10.425 0.980 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 7.245 2.010 7.575 2.980 ;
        RECT 8.195 2.010 8.525 2.980 ;
        RECT 7.245 1.840 8.525 2.010 ;
        RECT 8.285 1.170 8.525 1.840 ;
        RECT 7.265 0.920 8.615 1.170 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.115 2.255 0.445 2.980 ;
        RECT 0.645 2.425 0.815 3.245 ;
        RECT 0.985 2.630 2.005 2.960 ;
        RECT 0.985 2.255 1.155 2.630 ;
        RECT 2.210 2.460 2.540 2.755 ;
        RECT 0.115 2.085 1.155 2.255 ;
        RECT 1.325 2.290 2.540 2.460 ;
        RECT 0.115 1.950 0.445 2.085 ;
        RECT 1.325 1.915 1.495 2.290 ;
        RECT 3.170 2.085 3.500 3.245 ;
        RECT 3.670 2.255 4.000 2.755 ;
        RECT 4.170 2.425 4.570 3.245 ;
        RECT 4.740 2.255 5.070 2.755 ;
        RECT 3.670 2.085 5.070 2.255 ;
        RECT 5.240 2.230 5.570 2.755 ;
        RECT 6.795 2.290 7.045 3.245 ;
        RECT 5.240 2.120 6.425 2.230 ;
        RECT 7.775 2.180 8.025 3.245 ;
        RECT 5.240 2.060 7.075 2.120 ;
        RECT 6.255 1.950 7.075 2.060 ;
        RECT 1.005 1.745 1.495 1.915 ;
        RECT 1.005 1.090 1.175 1.745 ;
        RECT 2.005 1.180 2.275 1.780 ;
        RECT 6.905 1.670 7.075 1.950 ;
        RECT 8.725 1.820 8.975 3.245 ;
        RECT 9.675 2.160 9.925 3.245 ;
        RECT 10.625 1.820 10.875 3.245 ;
        RECT 3.005 1.260 3.740 1.575 ;
        RECT 3.005 1.180 3.215 1.260 ;
        RECT 4.930 1.220 5.260 1.550 ;
        RECT 4.930 1.090 5.255 1.220 ;
        RECT 5.430 1.180 5.745 1.550 ;
        RECT 6.905 1.340 8.105 1.670 ;
        RECT 6.905 1.090 7.075 1.340 ;
        RECT 0.115 0.750 0.445 1.075 ;
        RECT 1.005 1.010 1.835 1.090 ;
        RECT 3.385 1.010 5.255 1.090 ;
        RECT 5.915 1.010 7.075 1.090 ;
        RECT 1.005 0.920 5.255 1.010 ;
        RECT 1.665 0.840 3.555 0.920 ;
        RECT 0.115 0.670 1.495 0.750 ;
        RECT 0.115 0.580 1.965 0.670 ;
        RECT 0.115 0.350 0.445 0.580 ;
        RECT 0.625 0.085 1.155 0.410 ;
        RECT 1.325 0.350 1.965 0.580 ;
        RECT 2.135 0.350 2.465 0.840 ;
        RECT 3.175 0.085 3.505 0.670 ;
        RECT 3.725 0.580 4.915 0.750 ;
        RECT 3.725 0.350 3.975 0.580 ;
        RECT 4.155 0.085 4.485 0.410 ;
        RECT 4.665 0.350 4.915 0.580 ;
        RECT 5.085 0.425 5.255 0.920 ;
        RECT 5.425 0.920 7.075 1.010 ;
        RECT 8.965 1.320 9.955 1.650 ;
        RECT 5.425 0.840 6.085 0.920 ;
        RECT 5.425 0.595 5.675 0.840 ;
        RECT 8.965 0.750 9.135 1.320 ;
        RECT 6.255 0.580 9.135 0.750 ;
        RECT 6.255 0.425 6.425 0.580 ;
        RECT 5.085 0.255 6.425 0.425 ;
        RECT 6.755 0.085 7.085 0.410 ;
        RECT 7.775 0.085 8.105 0.410 ;
        RECT 8.795 0.085 9.125 0.410 ;
        RECT 9.735 0.085 9.985 0.810 ;
        RECT 10.595 0.085 10.925 1.170 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 2.075 1.210 2.245 1.380 ;
        RECT 3.035 1.210 3.205 1.380 ;
        RECT 5.435 1.210 5.605 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__fa_4

#--------EOF---------

MACRO sky130_fd_sc_hs__fah_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fah_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 12.820 1.470 13.490 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.723000 ;
    PORT
      LAYER li1 ;
        RECT 9.145 1.180 9.475 1.550 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.410 1.335 1.780 ;
    END
  END CI
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.290 1.600 1.430 ;
        RECT 4.375 1.395 5.315 1.605 ;
        RECT 4.375 1.305 6.220 1.395 ;
        RECT 4.375 1.295 6.755 1.305 ;
        RECT 3.165 1.290 6.755 1.295 ;
        RECT 0.005 1.240 6.755 1.290 ;
        RECT 8.195 1.240 10.085 1.320 ;
        RECT 0.005 1.140 12.355 1.240 ;
        RECT 0.005 0.245 13.915 1.140 ;
        RECT 0.000 0.000 13.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.940 14.110 3.520 ;
        RECT -0.190 1.660 4.165 1.940 ;
        RECT 5.525 1.660 14.110 1.940 ;
        RECT 5.525 1.605 12.450 1.660 ;
        RECT 9.485 1.530 12.450 1.605 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.920 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.674850 ;
    PORT
      LAYER li1 ;
        RECT 0.985 2.905 2.645 3.075 ;
        RECT 0.985 2.120 1.155 2.905 ;
        RECT 2.315 2.875 2.645 2.905 ;
        RECT 0.665 1.950 1.155 2.120 ;
        RECT 0.665 0.900 0.835 1.950 ;
        RECT 0.665 0.730 1.675 0.900 ;
        RECT 1.505 0.400 2.075 0.730 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.537600 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.540 0.445 2.980 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.920 3.415 ;
        RECT 0.645 2.290 0.815 3.245 ;
        RECT 2.935 2.965 3.290 3.245 ;
        RECT 3.460 2.905 7.000 3.075 ;
        RECT 3.460 2.795 3.630 2.905 ;
        RECT 1.325 2.705 1.675 2.735 ;
        RECT 2.815 2.705 3.630 2.795 ;
        RECT 1.325 2.625 3.630 2.705 ;
        RECT 1.325 2.535 2.985 2.625 ;
        RECT 1.325 1.950 1.675 2.535 ;
        RECT 4.205 2.455 4.535 2.735 ;
        RECT 3.155 2.365 4.535 2.455 ;
        RECT 1.505 1.240 1.675 1.950 ;
        RECT 1.130 1.070 1.675 1.240 ;
        RECT 1.845 2.285 4.535 2.365 ;
        RECT 1.845 2.195 3.325 2.285 ;
        RECT 1.845 1.070 2.175 2.195 ;
        RECT 3.495 2.025 4.000 2.115 ;
        RECT 4.205 2.100 4.535 2.285 ;
        RECT 4.705 2.730 6.125 2.905 ;
        RECT 3.005 1.855 4.000 2.025 ;
        RECT 2.500 1.410 2.830 1.635 ;
        RECT 3.005 1.580 3.445 1.855 ;
        RECT 4.705 1.765 4.875 2.730 ;
        RECT 6.330 2.490 6.660 2.640 ;
        RECT 4.170 1.685 4.875 1.765 ;
        RECT 2.500 1.240 3.105 1.410 ;
        RECT 1.845 0.900 2.765 1.070 ;
        RECT 0.620 0.085 0.950 0.560 ;
        RECT 2.255 0.085 2.425 0.730 ;
        RECT 2.595 0.425 2.765 0.900 ;
        RECT 2.935 0.765 3.105 1.240 ;
        RECT 3.275 1.185 3.445 1.580 ;
        RECT 3.670 1.595 4.875 1.685 ;
        RECT 5.045 2.320 6.660 2.490 ;
        RECT 3.670 1.435 4.340 1.595 ;
        RECT 5.045 1.425 5.215 2.320 ;
        RECT 6.330 2.290 6.660 2.320 ;
        RECT 4.880 1.265 5.215 1.425 ;
        RECT 5.405 1.705 5.635 2.150 ;
        RECT 6.830 2.120 7.000 2.905 ;
        RECT 6.055 1.950 7.000 2.120 ;
        RECT 7.170 1.950 7.500 2.925 ;
        RECT 5.405 1.375 5.885 1.705 ;
        RECT 3.275 0.935 3.605 1.185 ;
        RECT 3.775 1.095 5.215 1.265 ;
        RECT 6.055 1.205 6.225 1.950 ;
        RECT 3.775 0.765 3.945 1.095 ;
        RECT 5.385 1.035 6.225 1.205 ;
        RECT 6.395 1.550 6.595 1.780 ;
        RECT 6.845 1.550 7.075 1.780 ;
        RECT 5.385 0.935 5.715 1.035 ;
        RECT 2.935 0.595 3.945 0.765 ;
        RECT 4.115 0.765 5.045 0.925 ;
        RECT 5.885 0.765 6.215 0.865 ;
        RECT 4.115 0.755 6.215 0.765 ;
        RECT 4.115 0.425 4.285 0.755 ;
        RECT 4.875 0.595 6.215 0.755 ;
        RECT 6.395 0.670 6.565 1.550 ;
        RECT 6.845 1.380 7.065 1.550 ;
        RECT 6.735 0.710 7.065 1.380 ;
        RECT 7.330 1.130 7.500 1.950 ;
        RECT 7.670 1.765 8.000 3.245 ;
        RECT 8.170 2.905 11.740 3.075 ;
        RECT 8.170 1.880 8.610 2.905 ;
        RECT 8.780 2.565 10.815 2.735 ;
        RECT 8.780 1.880 9.110 2.565 ;
        RECT 8.170 1.210 8.340 1.880 ;
        RECT 9.280 1.805 10.475 2.395 ;
        RECT 8.510 1.380 8.975 1.710 ;
        RECT 7.235 0.790 7.565 1.130 ;
        RECT 8.170 0.960 8.635 1.210 ;
        RECT 8.805 0.790 8.975 1.380 ;
        RECT 9.645 0.960 9.975 1.805 ;
        RECT 10.145 1.220 10.475 1.550 ;
        RECT 10.145 0.790 10.315 1.220 ;
        RECT 10.645 1.050 10.815 2.565 ;
        RECT 7.235 0.620 10.315 0.790 ;
        RECT 2.595 0.255 4.285 0.425 ;
        RECT 4.455 0.425 4.705 0.585 ;
        RECT 7.235 0.425 7.565 0.620 ;
        RECT 10.485 0.595 10.815 1.050 ;
        RECT 10.985 1.780 11.155 2.735 ;
        RECT 10.985 1.550 11.215 1.780 ;
        RECT 4.455 0.255 7.565 0.425 ;
        RECT 7.745 0.085 8.075 0.450 ;
        RECT 8.895 0.425 9.385 0.450 ;
        RECT 10.985 0.425 11.155 1.550 ;
        RECT 11.385 1.130 11.740 2.905 ;
        RECT 11.950 2.330 12.290 3.245 ;
        RECT 11.950 2.110 12.220 2.330 ;
        RECT 12.520 2.160 12.850 2.980 ;
        RECT 12.390 1.970 12.850 2.160 ;
        RECT 13.050 1.970 13.300 3.245 ;
        RECT 13.470 1.970 13.830 2.980 ;
        RECT 12.390 1.940 12.650 1.970 ;
        RECT 8.895 0.255 11.155 0.425 ;
        RECT 11.405 0.350 11.740 1.130 ;
        RECT 11.910 1.720 12.650 1.940 ;
        RECT 11.910 0.960 12.080 1.720 ;
        RECT 12.250 1.300 12.580 1.550 ;
        RECT 13.660 1.300 13.830 1.970 ;
        RECT 12.250 1.130 13.830 1.300 ;
        RECT 11.910 0.790 12.805 0.960 ;
        RECT 11.915 0.085 12.245 0.620 ;
        RECT 12.475 0.350 12.805 0.790 ;
        RECT 12.975 0.085 13.305 0.960 ;
        RECT 13.475 0.350 13.830 1.130 ;
        RECT 0.000 -0.085 13.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 3.035 1.580 3.205 1.750 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 6.395 1.580 6.565 1.750 ;
        RECT 6.875 1.580 7.045 1.750 ;
        RECT 8.840 1.950 9.010 2.120 ;
        RECT 9.885 1.950 10.055 2.120 ;
        RECT 10.245 1.950 10.415 2.120 ;
        RECT 11.015 1.580 11.185 1.750 ;
        RECT 12.435 1.950 12.605 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
      LAYER met1 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 8.780 2.105 9.070 2.150 ;
        RECT 5.375 1.965 9.070 2.105 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 8.780 1.920 9.070 1.965 ;
        RECT 9.825 2.105 10.475 2.150 ;
        RECT 12.375 2.105 12.665 2.150 ;
        RECT 9.825 1.965 12.665 2.105 ;
        RECT 9.825 1.920 10.475 1.965 ;
        RECT 12.375 1.920 12.665 1.965 ;
        RECT 2.975 1.735 3.265 1.780 ;
        RECT 6.335 1.735 6.625 1.780 ;
        RECT 2.975 1.595 6.625 1.735 ;
        RECT 2.975 1.550 3.265 1.595 ;
        RECT 6.335 1.550 6.625 1.595 ;
        RECT 6.815 1.735 7.105 1.780 ;
        RECT 10.955 1.735 11.245 1.780 ;
        RECT 6.815 1.595 11.245 1.735 ;
        RECT 6.815 1.550 7.105 1.595 ;
        RECT 10.955 1.550 11.245 1.595 ;
  END
END sky130_fd_sc_hs__fah_1

#--------EOF---------

MACRO sky130_fd_sc_hs__fah_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fah_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.290 2.045 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.723000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.355 2.895 2.150 ;
        RECT 3.440 1.630 3.770 1.960 ;
        RECT 2.725 0.765 2.895 1.355 ;
        RECT 3.565 0.765 3.735 1.630 ;
        RECT 4.405 0.765 4.595 1.605 ;
        RECT 5.875 1.090 6.205 1.185 ;
        RECT 5.265 0.920 6.205 1.090 ;
        RECT 5.265 0.765 5.435 0.920 ;
        RECT 2.725 0.595 5.435 0.765 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 11.450 1.450 11.875 1.780 ;
    END
  END CI
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.265 1.240 5.745 1.295 ;
        RECT 0.080 0.940 5.745 1.240 ;
        RECT 6.670 1.165 7.580 1.240 ;
        RECT 9.475 1.165 10.025 1.295 ;
        RECT 11.975 1.165 14.395 1.240 ;
        RECT 6.670 0.940 14.395 1.165 ;
        RECT 0.080 0.245 14.395 0.940 ;
        RECT 0.000 0.000 14.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.400 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 12.585 1.550 12.920 2.200 ;
        RECT 12.585 0.350 12.835 1.550 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.561800 ;
    PORT
      LAYER li1 ;
        RECT 13.570 1.820 13.875 2.980 ;
        RECT 13.705 1.505 13.875 1.820 ;
        RECT 13.705 1.130 14.275 1.505 ;
        RECT 13.515 0.800 14.275 1.130 ;
        RECT 13.515 0.355 13.785 0.800 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.400 3.415 ;
        RECT 0.105 2.160 0.360 3.245 ;
        RECT 0.555 1.990 0.885 2.980 ;
        RECT 0.335 1.820 0.885 1.990 ;
        RECT 0.335 1.470 0.650 1.820 ;
        RECT 1.090 1.630 1.340 2.980 ;
        RECT 1.540 1.950 1.870 3.245 ;
        RECT 2.055 2.890 6.055 3.060 ;
        RECT 2.055 2.015 2.385 2.890 ;
        RECT 2.555 2.550 5.555 2.720 ;
        RECT 2.555 2.390 3.450 2.550 ;
        RECT 0.125 1.180 0.650 1.470 ;
        RECT 0.820 1.300 1.395 1.630 ;
        RECT 0.480 1.130 0.650 1.180 ;
        RECT 0.480 0.960 0.965 1.130 ;
        RECT 0.170 0.085 0.535 0.790 ;
        RECT 0.705 0.350 0.965 0.960 ;
        RECT 1.225 1.120 1.395 1.300 ;
        RECT 2.215 1.185 2.385 2.015 ;
        RECT 3.065 1.185 3.235 2.390 ;
        RECT 3.620 2.130 4.110 2.380 ;
        RECT 3.940 1.410 4.110 2.130 ;
        RECT 4.280 2.100 5.215 2.350 ;
        RECT 5.385 2.270 5.555 2.550 ;
        RECT 5.725 2.440 6.055 2.890 ;
        RECT 6.265 2.580 6.595 3.245 ;
        RECT 7.215 2.905 9.575 3.075 ;
        RECT 7.215 2.410 7.385 2.905 ;
        RECT 6.225 2.270 7.385 2.410 ;
        RECT 5.385 2.240 7.385 2.270 ;
        RECT 5.385 2.100 6.395 2.240 ;
        RECT 4.765 1.430 4.935 2.100 ;
        RECT 6.715 1.930 7.045 2.070 ;
        RECT 5.105 1.760 7.045 1.930 ;
        RECT 5.105 1.600 5.365 1.760 ;
        RECT 5.535 1.430 6.545 1.525 ;
        RECT 3.940 1.185 4.235 1.410 ;
        RECT 1.225 0.505 1.705 1.120 ;
        RECT 2.215 1.015 2.555 1.185 ;
        RECT 1.875 0.085 2.125 0.845 ;
        RECT 2.305 0.425 2.555 1.015 ;
        RECT 3.065 0.935 3.395 1.185 ;
        RECT 3.905 0.935 4.235 1.185 ;
        RECT 4.765 1.355 6.545 1.430 ;
        RECT 4.765 1.260 5.705 1.355 ;
        RECT 4.765 0.935 5.095 1.260 ;
        RECT 6.375 1.020 6.545 1.355 ;
        RECT 6.715 1.360 7.045 1.760 ;
        RECT 7.215 1.960 7.385 2.240 ;
        RECT 7.555 2.130 8.310 2.735 ;
        RECT 7.215 1.630 7.505 1.960 ;
        RECT 6.715 1.190 7.505 1.360 ;
        RECT 6.375 0.850 7.005 1.020 ;
        RECT 5.605 0.425 5.935 0.750 ;
        RECT 2.305 0.255 5.935 0.425 ;
        RECT 6.335 0.085 6.665 0.680 ;
        RECT 6.835 0.425 7.005 0.850 ;
        RECT 7.175 0.630 7.505 1.190 ;
        RECT 7.675 1.275 7.970 1.945 ;
        RECT 7.675 0.425 7.845 1.275 ;
        RECT 8.140 1.040 8.310 2.130 ;
        RECT 8.480 1.225 8.735 2.905 ;
        RECT 8.905 2.130 9.235 2.735 ;
        RECT 8.905 1.055 9.075 2.130 ;
        RECT 9.405 1.960 9.575 2.905 ;
        RECT 8.140 0.640 8.555 1.040 ;
        RECT 6.835 0.255 7.845 0.425 ;
        RECT 8.015 0.390 8.555 0.640 ;
        RECT 8.745 0.425 9.075 1.055 ;
        RECT 9.245 1.630 9.575 1.960 ;
        RECT 9.745 2.770 10.075 2.980 ;
        RECT 11.015 2.940 11.395 3.245 ;
        RECT 9.745 2.600 11.970 2.770 ;
        RECT 12.140 2.710 12.470 3.245 ;
        RECT 13.040 2.710 13.370 3.245 ;
        RECT 9.745 2.100 10.075 2.600 ;
        RECT 11.800 2.540 11.970 2.600 ;
        RECT 10.310 2.130 10.810 2.430 ;
        RECT 11.800 2.370 13.400 2.540 ;
        RECT 9.245 0.765 9.415 1.630 ;
        RECT 9.745 1.185 9.915 2.100 ;
        RECT 9.585 0.935 9.915 1.185 ;
        RECT 10.085 1.355 10.470 1.685 ;
        RECT 10.085 0.765 10.255 1.355 ;
        RECT 10.640 1.185 10.810 2.130 ;
        RECT 9.245 0.595 10.255 0.765 ;
        RECT 10.425 1.015 10.810 1.185 ;
        RECT 10.980 1.950 11.930 2.200 ;
        RECT 10.980 1.055 11.240 1.950 ;
        RECT 13.230 1.630 13.400 2.370 ;
        RECT 14.045 1.820 14.295 3.245 ;
        RECT 10.425 0.595 10.595 1.015 ;
        RECT 10.980 0.845 11.865 1.055 ;
        RECT 10.765 0.675 11.865 0.845 ;
        RECT 12.085 0.810 12.415 1.550 ;
        RECT 13.230 1.300 13.535 1.630 ;
        RECT 10.765 0.425 10.935 0.675 ;
        RECT 8.745 0.255 10.935 0.425 ;
        RECT 11.105 0.085 11.355 0.505 ;
        RECT 11.535 0.375 11.865 0.675 ;
        RECT 12.075 0.085 12.405 0.640 ;
        RECT 13.015 0.085 13.345 1.130 ;
        RECT 13.955 0.085 14.285 0.630 ;
        RECT 0.000 -0.085 14.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 0.155 1.210 0.325 1.380 ;
        RECT 3.995 1.210 4.165 1.380 ;
        RECT 8.315 0.840 8.485 1.010 ;
        RECT 12.155 0.840 12.325 1.010 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
      LAYER met1 ;
        RECT 0.095 1.365 0.385 1.410 ;
        RECT 3.935 1.365 4.225 1.410 ;
        RECT 0.095 1.225 4.225 1.365 ;
        RECT 0.095 1.180 0.385 1.225 ;
        RECT 3.935 1.180 4.225 1.225 ;
        RECT 8.255 0.995 8.545 1.040 ;
        RECT 12.095 0.995 12.385 1.040 ;
        RECT 8.255 0.855 12.385 0.995 ;
        RECT 8.255 0.810 8.545 0.855 ;
        RECT 12.095 0.810 12.385 0.855 ;
  END
END sky130_fd_sc_hs__fah_2

#--------EOF---------

MACRO sky130_fd_sc_hs__fah_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fah_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.510 1.095 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.723000 ;
    PORT
      LAYER li1 ;
        RECT 4.675 2.290 5.155 2.910 ;
        RECT 4.675 1.220 4.925 2.290 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 12.635 1.350 12.980 1.780 ;
    END
  END CI
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 15.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.090 1.340 4.485 1.420 ;
        RECT 7.265 1.395 8.190 1.505 ;
        RECT 1.425 1.240 4.485 1.340 ;
        RECT 6.360 1.375 8.190 1.395 ;
        RECT 6.360 1.370 9.405 1.375 ;
        RECT 6.360 1.280 15.355 1.370 ;
        RECT 5.785 1.240 15.355 1.280 ;
        RECT 1.425 1.140 15.355 1.240 ;
        RECT 0.005 0.245 15.355 1.140 ;
        RECT 0.000 0.000 15.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.715 15.550 3.520 ;
        RECT -0.190 1.660 7.055 1.715 ;
        RECT 8.400 1.660 15.550 1.715 ;
        RECT 1.415 1.630 7.055 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 15.360 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 9.890 1.850 11.395 2.100 ;
        RECT 10.960 1.260 11.395 1.850 ;
        RECT 10.960 1.180 11.785 1.260 ;
        RECT 10.475 1.010 11.785 1.180 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.097600 ;
    PORT
      LAYER li1 ;
        RECT 13.420 2.020 13.750 2.980 ;
        RECT 14.420 2.020 14.755 2.980 ;
        RECT 13.420 1.850 14.755 2.020 ;
        RECT 14.495 1.180 14.745 1.850 ;
        RECT 13.555 1.010 14.745 1.180 ;
        RECT 13.555 0.480 13.805 1.010 ;
        RECT 14.495 0.480 14.745 1.010 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 15.360 3.415 ;
        RECT 0.085 1.970 0.365 2.980 ;
        RECT 0.565 1.970 0.815 3.245 ;
        RECT 1.015 2.800 1.345 2.980 ;
        RECT 1.575 2.970 1.915 3.245 ;
        RECT 3.165 2.800 3.495 2.960 ;
        RECT 1.015 2.630 3.495 2.800 ;
        RECT 1.015 1.970 1.345 2.630 ;
        RECT 0.085 1.340 0.255 1.970 ;
        RECT 1.335 1.340 1.665 1.650 ;
        RECT 0.085 1.170 1.665 1.340 ;
        RECT 0.085 0.350 0.365 1.170 ;
        RECT 1.835 1.000 2.005 2.630 ;
        RECT 4.230 2.460 4.505 2.670 ;
        RECT 2.175 2.290 4.505 2.460 ;
        RECT 5.325 2.290 5.655 3.245 ;
        RECT 2.175 1.790 2.505 2.290 ;
        RECT 0.545 0.085 0.795 1.000 ;
        RECT 0.975 0.960 2.005 1.000 ;
        RECT 0.975 0.790 2.135 0.960 ;
        RECT 0.975 0.350 1.305 0.790 ;
        RECT 1.535 0.085 1.795 0.620 ;
        RECT 1.965 0.425 2.135 0.790 ;
        RECT 2.305 0.625 2.475 1.790 ;
        RECT 2.705 1.780 2.960 2.120 ;
        RECT 3.375 1.935 4.030 2.120 ;
        RECT 4.230 1.935 4.505 2.290 ;
        RECT 5.855 2.120 6.025 2.980 ;
        RECT 2.705 1.550 3.205 1.780 ;
        RECT 3.375 1.380 3.545 1.935 ;
        RECT 2.655 1.210 3.545 1.380 ;
        RECT 3.715 1.550 4.165 1.765 ;
        RECT 2.655 0.625 2.985 1.210 ;
        RECT 3.155 0.425 3.415 1.040 ;
        RECT 3.715 0.630 3.885 1.550 ;
        RECT 4.335 1.310 4.505 1.935 ;
        RECT 4.065 1.045 4.505 1.310 ;
        RECT 5.095 1.950 6.025 2.120 ;
        RECT 6.195 2.905 8.715 3.075 ;
        RECT 9.115 2.950 9.685 3.245 ;
        RECT 10.425 2.950 10.755 3.245 ;
        RECT 11.495 2.950 12.125 3.245 ;
        RECT 6.195 2.150 6.365 2.905 ;
        RECT 6.535 2.490 6.785 2.735 ;
        RECT 6.990 2.725 7.875 2.905 ;
        RECT 8.545 2.780 8.715 2.905 ;
        RECT 12.295 2.780 12.715 2.860 ;
        RECT 6.535 2.320 7.535 2.490 ;
        RECT 6.195 1.980 6.485 2.150 ;
        RECT 5.095 0.920 5.265 1.950 ;
        RECT 5.435 1.375 5.635 1.780 ;
        RECT 5.885 1.550 6.145 1.780 ;
        RECT 5.435 1.090 5.805 1.375 ;
        RECT 5.095 0.875 5.405 0.920 ;
        RECT 5.975 0.875 6.145 1.550 ;
        RECT 6.315 1.215 6.485 1.980 ;
        RECT 6.655 1.405 7.075 2.150 ;
        RECT 7.365 1.285 7.535 2.320 ;
        RECT 7.705 1.650 7.875 2.725 ;
        RECT 8.045 2.440 8.375 2.735 ;
        RECT 8.545 2.610 12.715 2.780 ;
        RECT 8.045 2.270 12.125 2.440 ;
        RECT 8.045 2.095 8.375 2.270 ;
        RECT 8.580 1.900 9.215 2.100 ;
        RECT 9.045 1.775 9.215 1.900 ;
        RECT 7.705 1.480 8.875 1.650 ;
        RECT 8.205 1.320 8.875 1.480 ;
        RECT 9.045 1.550 9.475 1.775 ;
        RECT 6.315 1.045 7.195 1.215 ;
        RECT 6.865 1.015 7.195 1.045 ;
        RECT 7.365 1.105 7.685 1.285 ;
        RECT 7.365 0.935 8.875 1.105 ;
        RECT 9.045 0.935 9.215 1.550 ;
        RECT 9.780 1.350 10.710 1.680 ;
        RECT 9.780 1.180 9.950 1.350 ;
        RECT 9.385 1.010 9.950 1.180 ;
        RECT 4.055 0.705 5.405 0.875 ;
        RECT 1.965 0.255 3.415 0.425 ;
        RECT 4.055 0.255 4.385 0.705 ;
        RECT 4.585 0.085 4.915 0.535 ;
        RECT 5.095 0.425 5.405 0.705 ;
        RECT 5.875 0.595 6.205 0.875 ;
        RECT 6.375 0.765 6.705 0.845 ;
        RECT 8.705 0.765 8.875 0.935 ;
        RECT 9.385 0.765 9.555 1.010 ;
        RECT 11.955 0.840 12.125 2.270 ;
        RECT 12.295 1.950 12.715 2.610 ;
        RECT 12.920 1.950 13.250 3.245 ;
        RECT 13.920 2.190 14.250 3.245 ;
        RECT 12.295 1.180 12.465 1.950 ;
        RECT 14.950 1.820 15.200 3.245 ;
        RECT 13.215 1.350 14.325 1.680 ;
        RECT 12.295 1.010 12.855 1.180 ;
        RECT 13.215 0.840 13.385 1.350 ;
        RECT 6.375 0.595 8.535 0.765 ;
        RECT 8.705 0.595 9.555 0.765 ;
        RECT 9.725 0.670 13.385 0.840 ;
        RECT 8.365 0.425 8.535 0.595 ;
        RECT 9.725 0.425 9.895 0.670 ;
        RECT 5.095 0.255 8.195 0.425 ;
        RECT 8.365 0.255 9.895 0.425 ;
        RECT 10.065 0.085 10.315 0.500 ;
        RECT 10.965 0.085 11.295 0.500 ;
        RECT 11.965 0.085 12.295 0.500 ;
        RECT 13.035 0.085 13.375 0.500 ;
        RECT 13.985 0.085 14.315 0.840 ;
        RECT 14.915 0.085 15.245 1.260 ;
        RECT 0.000 -0.085 15.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 3.515 1.950 3.685 2.120 ;
        RECT 3.035 1.580 3.205 1.750 ;
        RECT 3.995 1.580 4.165 1.750 ;
        RECT 5.435 1.580 5.605 1.750 ;
        RECT 5.915 1.580 6.085 1.750 ;
        RECT 6.875 1.950 7.045 2.120 ;
        RECT 9.275 1.580 9.445 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
      LAYER met1 ;
        RECT 3.455 2.105 3.745 2.150 ;
        RECT 6.815 2.105 7.105 2.150 ;
        RECT 3.455 1.965 7.105 2.105 ;
        RECT 3.455 1.920 3.745 1.965 ;
        RECT 6.815 1.920 7.105 1.965 ;
        RECT 2.975 1.735 3.265 1.780 ;
        RECT 3.935 1.735 4.225 1.780 ;
        RECT 5.375 1.735 5.665 1.780 ;
        RECT 2.975 1.595 5.665 1.735 ;
        RECT 2.975 1.550 3.265 1.595 ;
        RECT 3.935 1.550 4.225 1.595 ;
        RECT 5.375 1.550 5.665 1.595 ;
        RECT 5.855 1.735 6.145 1.780 ;
        RECT 9.215 1.735 9.505 1.780 ;
        RECT 5.855 1.595 9.505 1.735 ;
        RECT 5.855 1.550 6.145 1.595 ;
        RECT 9.215 1.550 9.505 1.595 ;
  END
END sky130_fd_sc_hs__fah_4

#--------EOF---------

MACRO sky130_fd_sc_hs__fahcin_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fahcin_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.350 0.835 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.723000 ;
    PORT
      LAYER li1 ;
        RECT 4.875 1.180 5.205 1.585 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.525000 ;
    PORT
      LAYER li1 ;
        RECT 8.705 1.155 9.035 1.485 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.015 1.370 11.345 1.450 ;
        RECT 3.155 1.275 4.815 1.365 ;
        RECT 0.010 1.140 1.900 1.240 ;
        RECT 3.155 1.175 5.815 1.275 ;
        RECT 9.015 1.175 12.955 1.370 ;
        RECT 3.155 1.140 12.955 1.175 ;
        RECT 0.010 0.245 12.955 1.140 ;
        RECT 0.000 0.000 12.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.150 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.960 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.959800 ;
    PORT
      LAYER li1 ;
        RECT 6.820 2.335 7.615 2.665 ;
        RECT 6.900 1.310 7.070 2.335 ;
        RECT 6.640 0.985 7.070 1.310 ;
        RECT 6.640 0.440 8.035 0.985 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 12.595 0.840 12.845 2.980 ;
        RECT 12.515 0.440 12.845 0.840 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.120 1.180 0.375 2.980 ;
        RECT 0.575 1.950 0.825 3.245 ;
        RECT 1.005 2.905 3.935 3.075 ;
        RECT 1.005 1.630 1.175 2.905 ;
        RECT 1.345 2.565 2.980 2.735 ;
        RECT 1.345 1.820 1.835 2.565 ;
        RECT 2.045 2.070 2.485 2.395 ;
        RECT 2.045 1.890 2.415 2.070 ;
        RECT 2.655 2.045 2.980 2.565 ;
        RECT 1.005 1.300 1.445 1.630 ;
        RECT 1.005 1.180 1.290 1.300 ;
        RECT 0.120 1.010 1.290 1.180 ;
        RECT 1.615 1.020 1.835 1.820 ;
        RECT 0.120 0.350 0.450 1.010 ;
        RECT 0.620 0.085 0.950 0.840 ;
        RECT 1.120 0.425 1.290 1.010 ;
        RECT 1.475 0.615 1.835 1.020 ;
        RECT 2.165 0.615 2.415 1.890 ;
        RECT 2.810 1.090 2.980 2.045 ;
        RECT 3.185 2.050 3.515 2.735 ;
        RECT 3.685 2.250 3.935 2.905 ;
        RECT 4.105 2.905 5.045 3.075 ;
        RECT 4.105 2.050 4.275 2.905 ;
        RECT 3.185 1.880 4.275 2.050 ;
        RECT 3.185 1.875 3.515 1.880 ;
        RECT 4.445 1.875 4.705 2.735 ;
        RECT 4.875 2.560 5.045 2.905 ;
        RECT 5.405 2.730 5.765 3.245 ;
        RECT 6.150 2.905 8.715 3.075 ;
        RECT 6.150 2.560 6.650 2.905 ;
        RECT 4.875 2.390 6.650 2.560 ;
        RECT 2.810 0.920 3.175 1.090 ;
        RECT 2.585 0.425 2.835 0.750 ;
        RECT 1.120 0.255 2.835 0.425 ;
        RECT 3.005 0.425 3.175 0.920 ;
        RECT 3.345 0.595 3.515 1.875 ;
        RECT 3.685 1.550 3.990 1.710 ;
        RECT 3.685 1.380 4.285 1.550 ;
        RECT 3.695 0.425 3.945 1.125 ;
        RECT 3.005 0.255 3.945 0.425 ;
        RECT 4.115 0.425 4.285 1.380 ;
        RECT 4.455 0.670 4.705 1.875 ;
        RECT 4.955 1.990 5.285 2.220 ;
        RECT 4.955 1.820 5.800 1.990 ;
        RECT 5.970 1.820 6.310 2.220 ;
        RECT 5.630 1.585 5.800 1.820 ;
        RECT 5.630 1.255 5.970 1.585 ;
        RECT 5.630 1.010 5.800 1.255 ;
        RECT 4.965 0.840 5.800 1.010 ;
        RECT 6.140 1.065 6.310 1.820 ;
        RECT 6.480 1.840 6.650 2.390 ;
        RECT 6.480 1.510 6.730 1.840 ;
        RECT 7.240 1.170 7.555 2.150 ;
        RECT 7.785 1.485 7.955 2.905 ;
        RECT 8.125 1.820 8.375 2.735 ;
        RECT 7.745 1.155 8.035 1.485 ;
        RECT 8.205 1.065 8.375 1.820 ;
        RECT 8.545 1.825 8.715 2.905 ;
        RECT 8.885 1.995 9.055 3.245 ;
        RECT 9.255 2.905 11.975 3.075 ;
        RECT 9.255 1.995 9.725 2.905 ;
        RECT 10.800 2.740 11.155 2.905 ;
        RECT 8.545 1.655 9.385 1.825 ;
        RECT 4.965 0.425 5.295 0.840 ;
        RECT 4.115 0.255 5.295 0.425 ;
        RECT 5.465 0.085 5.970 0.635 ;
        RECT 6.140 0.385 6.470 1.065 ;
        RECT 8.205 0.385 8.535 1.065 ;
        RECT 8.705 0.085 9.045 0.985 ;
        RECT 9.215 0.570 9.385 1.655 ;
        RECT 9.555 1.340 9.725 1.995 ;
        RECT 9.895 2.570 10.065 2.735 ;
        RECT 11.385 2.570 11.635 2.735 ;
        RECT 9.895 2.400 11.635 2.570 ;
        RECT 9.895 1.900 10.065 2.400 ;
        RECT 9.555 0.740 9.885 1.340 ;
        RECT 10.265 1.260 10.515 2.230 ;
        RECT 10.685 1.430 11.015 2.150 ;
        RECT 11.195 1.850 11.635 2.400 ;
        RECT 10.070 0.740 10.915 1.260 ;
        RECT 11.195 1.250 11.365 1.850 ;
        RECT 11.805 1.680 11.975 2.905 ;
        RECT 12.145 1.850 12.395 3.245 ;
        RECT 11.535 1.350 11.975 1.680 ;
        RECT 9.215 0.255 10.575 0.570 ;
        RECT 10.745 0.490 10.915 0.740 ;
        RECT 11.085 1.220 11.365 1.250 ;
        RECT 11.085 0.660 11.415 1.220 ;
        RECT 12.145 1.180 12.425 1.680 ;
        RECT 11.585 1.010 12.425 1.180 ;
        RECT 11.585 0.490 11.755 1.010 ;
        RECT 10.745 0.320 11.755 0.490 ;
        RECT 11.925 0.085 12.345 0.810 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 2.075 1.950 2.245 2.120 ;
        RECT 4.475 1.950 4.645 2.120 ;
        RECT 7.355 1.950 7.525 2.120 ;
        RECT 10.715 1.950 10.885 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
      LAYER met1 ;
        RECT 2.015 2.105 2.305 2.150 ;
        RECT 4.415 2.105 4.705 2.150 ;
        RECT 7.295 2.105 7.585 2.150 ;
        RECT 10.655 2.105 10.945 2.150 ;
        RECT 2.015 1.965 10.945 2.105 ;
        RECT 2.015 1.920 2.305 1.965 ;
        RECT 4.415 1.920 4.705 1.965 ;
        RECT 7.295 1.920 7.585 1.965 ;
        RECT 10.655 1.920 10.945 1.965 ;
  END
END sky130_fd_sc_hs__fahcin_1

#--------EOF---------

MACRO sky130_fd_sc_hs__fahcon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fahcon_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.350 0.805 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.969000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.180 5.060 1.550 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.525000 ;
    PORT
      LAYER li1 ;
        RECT 7.675 1.180 8.005 1.550 ;
    END
  END CI
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.520 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.815 1.370 3.920 1.435 ;
        RECT 0.005 1.240 3.920 1.370 ;
        RECT 0.005 1.140 5.265 1.240 ;
        RECT 7.680 1.140 11.515 1.240 ;
        RECT 0.005 0.245 11.515 1.140 ;
        RECT 0.000 0.000 11.520 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.710 3.520 ;
        RECT 1.250 1.645 5.035 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.520 3.575 ;
    END
  END VPWR
  PIN COUT_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.782600 ;
    PORT
      LAYER li1 ;
        RECT 5.790 2.255 6.120 2.965 ;
        RECT 5.790 2.085 6.175 2.255 ;
        RECT 6.005 1.380 6.175 2.085 ;
        RECT 6.005 1.210 6.650 1.380 ;
        RECT 6.320 0.350 6.650 1.210 ;
    END
  END COUT_N
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 11.075 1.820 11.435 2.980 ;
        RECT 11.265 1.130 11.435 1.820 ;
        RECT 11.155 0.350 11.435 1.130 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.085 1.950 0.485 2.980 ;
        RECT 0.655 1.950 0.985 3.245 ;
        RECT 1.190 2.905 3.810 3.075 ;
        RECT 0.085 1.180 0.255 1.950 ;
        RECT 1.190 1.850 1.520 2.905 ;
        RECT 0.975 1.180 1.180 1.680 ;
        RECT 1.350 1.490 1.520 1.850 ;
        RECT 1.690 2.565 3.260 2.735 ;
        RECT 1.690 1.830 1.860 2.565 ;
        RECT 2.030 2.225 3.275 2.395 ;
        RECT 2.030 2.000 2.200 2.225 ;
        RECT 1.690 1.660 2.095 1.830 ;
        RECT 2.400 1.805 2.775 2.055 ;
        RECT 1.350 1.320 1.745 1.490 ;
        RECT 0.085 1.150 1.180 1.180 ;
        RECT 0.085 0.980 1.245 1.150 ;
        RECT 0.085 0.480 0.365 0.980 ;
        RECT 0.545 0.480 0.905 0.810 ;
        RECT 0.545 0.085 0.715 0.480 ;
        RECT 1.075 0.425 1.245 0.980 ;
        RECT 1.415 0.595 1.745 1.320 ;
        RECT 1.925 1.325 2.095 1.660 ;
        RECT 1.925 0.595 2.275 1.325 ;
        RECT 2.445 0.725 2.775 1.805 ;
        RECT 2.945 0.725 3.275 2.225 ;
        RECT 2.445 0.425 2.615 0.725 ;
        RECT 3.460 0.645 3.810 2.905 ;
        RECT 4.040 1.805 4.375 2.965 ;
        RECT 4.545 1.805 4.875 3.245 ;
        RECT 5.100 1.975 5.430 2.965 ;
        RECT 6.345 2.085 7.475 2.970 ;
        RECT 4.040 1.010 4.210 1.805 ;
        RECT 5.230 1.305 5.400 1.975 ;
        RECT 5.570 1.475 5.835 1.805 ;
        RECT 6.345 1.550 6.610 1.880 ;
        RECT 5.230 1.135 5.495 1.305 ;
        RECT 1.075 0.255 2.615 0.425 ;
        RECT 2.785 0.425 3.115 0.555 ;
        RECT 4.040 0.425 4.735 1.010 ;
        RECT 2.785 0.255 4.735 0.425 ;
        RECT 4.905 0.085 5.155 0.965 ;
        RECT 5.325 0.640 5.495 1.135 ;
        RECT 5.665 1.040 5.835 1.475 ;
        RECT 6.820 1.130 7.135 1.800 ;
        RECT 5.665 0.810 6.115 1.040 ;
        RECT 6.820 0.810 7.075 1.130 ;
        RECT 7.305 0.960 7.475 2.085 ;
        RECT 7.645 1.940 7.815 3.245 ;
        RECT 8.015 2.490 8.345 2.980 ;
        RECT 8.575 2.870 10.455 3.040 ;
        RECT 8.575 2.660 8.905 2.870 ;
        RECT 9.560 2.490 10.030 2.700 ;
        RECT 8.015 2.320 10.030 2.490 ;
        RECT 8.015 1.820 8.345 2.320 ;
        RECT 8.175 1.130 8.345 1.820 ;
        RECT 9.135 1.820 9.360 2.150 ;
        RECT 9.560 1.820 10.030 2.320 ;
        RECT 8.515 1.550 8.965 1.780 ;
        RECT 8.515 1.300 8.765 1.550 ;
        RECT 9.135 1.380 9.305 1.820 ;
        RECT 9.860 1.590 10.030 1.820 ;
        RECT 10.200 1.930 10.455 2.870 ;
        RECT 10.650 2.100 10.900 3.245 ;
        RECT 10.200 1.760 10.625 1.930 ;
        RECT 8.935 1.210 9.305 1.380 ;
        RECT 9.475 1.260 9.690 1.590 ;
        RECT 9.860 1.260 10.285 1.590 ;
        RECT 8.935 1.130 9.105 1.210 ;
        RECT 5.325 0.390 6.150 0.640 ;
        RECT 7.245 0.350 7.575 0.960 ;
        RECT 7.745 0.085 7.995 1.010 ;
        RECT 8.175 0.350 8.515 1.130 ;
        RECT 8.775 0.425 9.105 1.130 ;
        RECT 9.475 1.040 9.645 1.260 ;
        RECT 10.455 1.090 10.625 1.760 ;
        RECT 9.275 0.810 9.645 1.040 ;
        RECT 9.815 0.920 10.625 1.090 ;
        RECT 10.810 1.300 11.095 1.630 ;
        RECT 9.815 0.595 9.985 0.920 ;
        RECT 10.810 0.750 10.980 1.300 ;
        RECT 10.155 0.580 10.980 0.750 ;
        RECT 10.155 0.425 10.325 0.580 ;
        RECT 8.775 0.255 10.325 0.425 ;
        RECT 10.495 0.085 10.895 0.410 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 2.075 0.840 2.245 1.010 ;
        RECT 3.035 1.580 3.205 1.750 ;
        RECT 6.395 1.580 6.565 1.750 ;
        RECT 5.915 0.840 6.085 1.010 ;
        RECT 6.875 0.840 7.045 1.010 ;
        RECT 8.795 1.580 8.965 1.750 ;
        RECT 9.275 0.840 9.445 1.010 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
      LAYER met1 ;
        RECT 2.975 1.735 3.265 1.780 ;
        RECT 6.335 1.735 6.625 1.780 ;
        RECT 8.735 1.735 9.025 1.780 ;
        RECT 2.975 1.595 9.025 1.735 ;
        RECT 2.975 1.550 3.265 1.595 ;
        RECT 6.335 1.550 6.625 1.595 ;
        RECT 8.735 1.550 9.025 1.595 ;
        RECT 2.015 0.995 2.305 1.040 ;
        RECT 5.855 0.995 6.145 1.040 ;
        RECT 6.815 0.995 7.105 1.040 ;
        RECT 9.215 0.995 9.505 1.040 ;
        RECT 2.015 0.855 9.505 0.995 ;
        RECT 2.015 0.810 2.305 0.855 ;
        RECT 5.855 0.810 6.145 0.855 ;
        RECT 6.815 0.810 7.105 0.855 ;
        RECT 9.215 0.810 9.505 0.855 ;
  END
END sky130_fd_sc_hs__fahcon_1

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.480 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.000 0.480 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 0.670 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.480 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.480 3.415 ;
        RECT 0.000 -0.085 0.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
  END
END sky130_fd_sc_hs__fill_1

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.000 0.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.150 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.960 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.960 3.415 ;
        RECT 0.000 -0.085 0.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
  END
END sky130_fd_sc_hs__fill_2

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__fill_4

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__fill_8

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_diode_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 0.955 1.240 ;
        RECT 0.000 0.000 0.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.150 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.960 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.960 3.415 ;
        RECT 0.135 2.750 0.825 3.245 ;
        RECT 0.135 0.085 0.825 0.580 ;
        RECT 0.000 -0.085 0.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
  END
END sky130_fd_sc_hs__fill_diode_2

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_diode_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_diode_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 1.915 1.240 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.135 2.750 1.785 3.245 ;
        RECT 0.135 0.085 1.785 0.580 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__fill_diode_4

#--------EOF---------

MACRO sky130_fd_sc_hs__fill_diode_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hs__fill_diode_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.135 2.750 3.705 3.245 ;
        RECT 0.135 0.085 3.705 0.580 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__fill_diode_8

#--------EOF---------

MACRO sky130_fd_sc_hs__ha_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ha_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.468000 ;
    PORT
      LAYER li1 ;
        RECT 2.450 0.255 2.780 0.670 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.468000 ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.550 3.300 1.800 ;
        RECT 1.765 1.470 2.095 1.550 ;
        RECT 2.970 1.470 3.300 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.955 1.420 2.900 1.465 ;
        RECT 0.960 1.365 2.900 1.420 ;
        RECT 0.960 1.240 4.750 1.365 ;
        RECT 0.005 0.245 4.750 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.780 4.990 3.520 ;
        RECT -0.190 1.660 1.745 1.780 ;
        RECT 3.110 1.660 4.990 1.780 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 4.310 1.850 4.715 2.980 ;
        RECT 4.545 1.180 4.715 1.850 ;
        RECT 4.310 0.475 4.715 1.180 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.820 0.445 2.980 ;
        RECT 0.115 1.130 0.355 1.820 ;
        RECT 0.115 0.350 0.445 1.130 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.615 2.650 1.205 3.245 ;
        RECT 1.410 2.480 1.740 2.800 ;
        RECT 0.685 2.310 1.740 2.480 ;
        RECT 2.485 2.310 3.190 3.245 ;
        RECT 0.685 1.630 0.855 2.310 ;
        RECT 3.360 2.140 3.640 2.980 ;
        RECT 0.525 1.300 0.855 1.630 ;
        RECT 1.195 1.970 3.640 2.140 ;
        RECT 3.810 2.100 4.140 3.245 ;
        RECT 1.195 1.470 1.525 1.970 ;
        RECT 3.470 1.680 3.640 1.970 ;
        RECT 2.460 1.300 2.790 1.355 ;
        RECT 0.685 1.130 1.400 1.300 ;
        RECT 1.070 0.910 1.400 1.130 ;
        RECT 1.580 1.130 2.790 1.300 ;
        RECT 3.470 1.350 4.375 1.680 ;
        RECT 3.470 1.255 3.640 1.350 ;
        RECT 0.625 0.085 0.875 0.795 ;
        RECT 1.580 0.630 1.750 1.130 ;
        RECT 1.930 0.085 2.280 0.960 ;
        RECT 2.460 0.840 2.790 1.130 ;
        RECT 3.020 1.085 3.640 1.255 ;
        RECT 3.020 0.575 3.350 1.085 ;
        RECT 3.810 0.085 4.140 1.180 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__ha_1

#--------EOF---------

MACRO sky130_fd_sc_hs__ha_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ha_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.450 1.390 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 2.320 2.120 2.520 ;
        RECT 0.125 1.630 0.295 2.320 ;
        RECT 0.125 1.300 0.550 1.630 ;
        RECT 1.790 1.450 2.120 2.320 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 4.865 1.820 5.195 2.170 ;
        RECT 4.885 1.130 5.055 1.820 ;
        RECT 4.885 0.350 5.215 1.130 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580200 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.820 4.675 2.170 ;
        RECT 4.505 1.050 4.675 1.820 ;
        RECT 3.975 0.880 4.675 1.050 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 2.690 0.445 3.245 ;
        RECT 1.015 2.690 1.400 3.245 ;
        RECT 3.080 2.680 3.845 3.245 ;
        RECT 4.415 2.680 4.745 3.245 ;
        RECT 5.315 2.680 5.645 3.245 ;
        RECT 2.290 2.340 5.555 2.510 ;
        RECT 0.565 1.980 0.895 2.150 ;
        RECT 0.720 1.280 0.890 1.980 ;
        RECT 2.290 1.610 2.460 2.340 ;
        RECT 2.630 1.920 3.490 2.170 ;
        RECT 2.290 1.280 3.035 1.610 ;
        RECT 3.320 1.550 3.490 1.920 ;
        RECT 5.385 1.630 5.555 2.340 ;
        RECT 0.720 1.130 2.460 1.280 ;
        RECT 0.115 1.110 2.460 1.130 ;
        RECT 3.320 1.220 4.330 1.550 ;
        RECT 5.225 1.300 5.555 1.630 ;
        RECT 3.320 1.110 3.490 1.220 ;
        RECT 0.115 0.960 0.890 1.110 ;
        RECT 0.115 0.350 0.445 0.960 ;
        RECT 2.635 0.940 3.490 1.110 ;
        RECT 1.365 0.770 2.465 0.940 ;
        RECT 0.935 0.085 1.265 0.600 ;
        RECT 1.795 0.085 2.125 0.600 ;
        RECT 2.295 0.425 2.465 0.770 ;
        RECT 2.635 0.595 2.805 0.940 ;
        RECT 2.985 0.425 3.315 0.770 ;
        RECT 2.295 0.255 3.315 0.425 ;
        RECT 3.545 0.085 3.875 0.710 ;
        RECT 4.455 0.085 4.705 0.710 ;
        RECT 5.395 0.085 5.645 1.130 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__ha_2

#--------EOF---------

MACRO sky130_fd_sc_hs__ha_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__ha_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.936000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.455 1.315 1.785 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.936000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.455 2.275 1.785 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.365 3.260 1.395 ;
        RECT 0.005 1.240 5.810 1.365 ;
        RECT 0.005 0.245 9.995 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
        RECT 3.545 1.585 4.805 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.265600 ;
    PORT
      LAYER li1 ;
        RECT 6.220 1.820 7.555 2.150 ;
        RECT 7.210 1.130 7.555 1.820 ;
        RECT 6.350 0.880 7.555 1.130 ;
        RECT 6.350 0.350 6.600 0.880 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.470100 ;
    PORT
      LAYER met1 ;
        RECT 8.735 2.105 9.025 2.150 ;
        RECT 9.695 2.105 9.985 2.150 ;
        RECT 8.735 1.965 9.985 2.105 ;
        RECT 8.735 1.920 9.025 1.965 ;
        RECT 9.695 1.920 9.985 1.965 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.105 2.125 0.385 2.965 ;
        RECT 0.555 2.295 0.805 3.245 ;
        RECT 1.005 2.905 2.235 3.075 ;
        RECT 1.005 2.125 1.255 2.905 ;
        RECT 0.105 1.955 1.255 2.125 ;
        RECT 1.455 2.125 1.735 2.735 ;
        RECT 1.905 2.295 2.235 2.905 ;
        RECT 2.475 2.405 2.805 3.245 ;
        RECT 3.375 2.505 3.705 3.245 ;
        RECT 4.430 2.660 4.760 3.245 ;
        RECT 5.490 2.660 5.945 3.245 ;
        RECT 6.675 2.660 7.005 3.245 ;
        RECT 7.575 2.660 7.905 3.245 ;
        RECT 3.900 2.335 7.895 2.490 ;
        RECT 3.085 2.320 7.895 2.335 ;
        RECT 3.085 2.235 4.070 2.320 ;
        RECT 2.925 2.165 4.070 2.235 ;
        RECT 2.925 2.125 3.255 2.165 ;
        RECT 1.455 1.955 3.255 2.125 ;
        RECT 4.955 1.995 6.050 2.150 ;
        RECT 2.500 1.905 3.255 1.955 ;
        RECT 2.500 1.285 2.670 1.905 ;
        RECT 3.900 1.820 6.050 1.995 ;
        RECT 3.900 1.745 4.230 1.820 ;
        RECT 3.900 1.735 4.070 1.745 ;
        RECT 3.075 1.575 4.070 1.735 ;
        RECT 5.880 1.650 6.050 1.820 ;
        RECT 7.725 1.650 7.895 2.320 ;
        RECT 8.075 2.150 8.305 2.980 ;
        RECT 8.475 2.320 8.805 3.245 ;
        RECT 9.075 2.150 9.405 2.980 ;
        RECT 9.635 2.320 9.965 3.245 ;
        RECT 8.075 1.820 9.995 2.150 ;
        RECT 3.075 1.405 4.280 1.575 ;
        RECT 0.115 1.115 2.170 1.285 ;
        RECT 0.115 0.605 0.365 1.115 ;
        RECT 0.545 0.085 0.795 0.945 ;
        RECT 0.980 0.605 1.230 1.115 ;
        RECT 1.410 0.085 1.660 0.945 ;
        RECT 1.840 0.435 2.170 1.115 ;
        RECT 2.340 0.605 2.670 1.285 ;
        RECT 2.840 0.435 3.170 1.235 ;
        RECT 1.840 0.265 3.170 0.435 ;
        RECT 3.520 0.485 3.780 1.235 ;
        RECT 3.950 0.655 4.280 1.405 ;
        RECT 4.450 1.425 5.710 1.595 ;
        RECT 4.450 0.485 4.780 1.425 ;
        RECT 3.520 0.315 4.780 0.485 ;
        RECT 4.950 0.085 5.280 1.255 ;
        RECT 5.460 0.575 5.710 1.425 ;
        RECT 5.880 1.320 6.955 1.650 ;
        RECT 7.725 1.320 9.645 1.650 ;
        RECT 9.825 1.150 9.995 1.820 ;
        RECT 5.920 0.085 6.170 1.130 ;
        RECT 8.150 0.980 9.995 1.150 ;
        RECT 6.780 0.085 7.110 0.710 ;
        RECT 7.640 0.085 7.970 0.710 ;
        RECT 8.150 0.350 8.400 0.980 ;
        RECT 8.570 0.085 8.900 0.810 ;
        RECT 9.070 0.350 9.400 0.980 ;
        RECT 9.580 0.085 9.885 0.810 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 8.795 1.950 8.965 2.120 ;
        RECT 9.755 1.950 9.925 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__ha_4

#--------EOF---------

MACRO sky130_fd_sc_hs__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.815 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.375 0.245 1.425 1.240 ;
        RECT 0.000 0.000 1.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.440 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.350 1.315 2.980 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.440 3.415 ;
        RECT 0.485 1.950 0.815 3.245 ;
        RECT 0.485 0.085 0.815 1.130 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
  END
END sky130_fd_sc_hs__inv_1

#--------EOF---------

MACRO sky130_fd_sc_hs__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 1.430 1.240 ;
        RECT 0.000 0.000 1.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.440 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.130 0.890 2.980 ;
        RECT 0.560 0.350 0.890 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.440 3.415 ;
        RECT 0.105 1.950 0.435 3.245 ;
        RECT 1.085 1.820 1.335 3.245 ;
        RECT 0.130 0.085 0.380 1.130 ;
        RECT 1.070 0.085 1.320 1.130 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
  END
END sky130_fd_sc_hs__inv_2

#--------EOF---------

MACRO sky130_fd_sc_hs__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.800 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 2.120 0.930 2.980 ;
        RECT 1.500 2.120 1.830 2.980 ;
        RECT 0.600 1.950 2.275 2.120 ;
        RECT 2.045 1.180 2.275 1.950 ;
        RECT 0.615 1.010 2.275 1.180 ;
        RECT 0.615 0.350 0.865 1.010 ;
        RECT 1.605 0.350 1.775 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.150 1.950 0.400 3.245 ;
        RECT 1.130 2.290 1.300 3.245 ;
        RECT 2.030 2.290 2.280 3.245 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 1.045 0.085 1.375 0.840 ;
        RECT 1.955 0.085 2.285 0.840 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__inv_4

#--------EOF---------

MACRO sky130_fd_sc_hs__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.232000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.350 2.250 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 4.225 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.172800 ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.120 0.815 2.980 ;
        RECT 1.515 2.120 1.845 2.980 ;
        RECT 2.495 2.120 2.665 2.980 ;
        RECT 0.565 1.950 2.665 2.120 ;
        RECT 2.495 1.620 2.665 1.950 ;
        RECT 3.365 1.620 3.695 2.980 ;
        RECT 2.495 1.310 4.195 1.620 ;
        RECT 2.420 1.180 4.195 1.310 ;
        RECT 0.560 1.140 4.195 1.180 ;
        RECT 0.560 1.010 2.680 1.140 ;
        RECT 0.560 0.350 0.810 1.010 ;
        RECT 1.500 0.350 1.670 1.010 ;
        RECT 2.350 0.350 2.680 1.010 ;
        RECT 3.350 0.350 3.610 1.140 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.015 2.290 1.345 3.245 ;
        RECT 2.045 2.290 2.295 3.245 ;
        RECT 2.865 1.820 3.195 3.245 ;
        RECT 3.865 1.820 4.195 3.245 ;
        RECT 0.130 0.085 0.380 1.130 ;
        RECT 0.990 0.085 1.320 0.840 ;
        RECT 1.850 0.085 2.180 0.840 ;
        RECT 2.850 0.085 3.180 0.970 ;
        RECT 3.780 0.085 4.110 0.970 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__inv_8

#--------EOF---------

MACRO sky130_fd_sc_hs__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.464000 ;
    PORT
      LAYER met1 ;
        RECT 1.085 1.550 7.070 1.780 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.095 0.245 8.065 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.379200 ;
    PORT
      LAYER met1 ;
        RECT 0.585 1.920 7.575 2.150 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 0.565 1.330 0.885 2.995 ;
        RECT 1.055 1.940 1.345 3.245 ;
        RECT 1.515 1.940 1.845 2.980 ;
        RECT 2.045 1.940 2.295 3.245 ;
        RECT 2.465 1.940 2.795 2.980 ;
        RECT 2.995 1.940 3.245 3.245 ;
        RECT 1.070 1.350 1.380 1.770 ;
        RECT 0.615 1.130 0.885 1.330 ;
        RECT 0.185 0.085 0.445 1.130 ;
        RECT 0.615 0.350 0.945 1.130 ;
        RECT 1.115 0.085 1.375 1.130 ;
        RECT 1.555 0.350 1.845 1.940 ;
        RECT 2.020 1.350 2.310 1.770 ;
        RECT 2.025 0.085 2.305 1.130 ;
        RECT 2.485 0.350 2.795 1.940 ;
        RECT 2.970 1.350 3.245 1.770 ;
        RECT 2.975 0.085 3.245 1.130 ;
        RECT 3.415 0.350 3.710 2.980 ;
        RECT 3.915 1.940 4.150 3.245 ;
        RECT 4.340 1.940 4.630 2.980 ;
        RECT 4.810 1.940 5.095 3.245 ;
        RECT 3.885 1.350 4.165 1.770 ;
        RECT 3.890 0.085 4.150 1.130 ;
        RECT 4.340 0.350 4.595 1.940 ;
        RECT 4.770 1.350 5.085 1.770 ;
        RECT 5.265 1.285 5.580 2.980 ;
        RECT 5.765 1.940 6.095 3.245 ;
        RECT 5.755 1.350 6.090 1.770 ;
        RECT 6.265 1.285 6.595 2.980 ;
        RECT 6.765 1.940 7.095 3.245 ;
        RECT 6.770 1.350 7.090 1.770 ;
        RECT 5.265 1.180 5.525 1.285 ;
        RECT 6.265 1.180 6.525 1.285 ;
        RECT 4.765 0.085 5.025 1.130 ;
        RECT 5.215 0.350 5.525 1.180 ;
        RECT 5.705 0.085 6.025 1.130 ;
        RECT 6.195 0.350 6.525 1.180 ;
        RECT 7.265 1.130 7.545 2.980 ;
        RECT 7.735 1.820 8.045 3.245 ;
        RECT 6.705 0.085 7.045 1.130 ;
        RECT 7.215 0.350 7.545 1.130 ;
        RECT 7.715 0.085 8.045 1.130 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.645 1.950 0.815 2.120 ;
        RECT 1.595 1.950 1.765 2.120 ;
        RECT 2.545 1.950 2.715 2.120 ;
        RECT 3.495 1.950 3.665 2.120 ;
        RECT 1.145 1.580 1.315 1.750 ;
        RECT 2.085 1.580 2.255 1.750 ;
        RECT 3.025 1.580 3.195 1.750 ;
        RECT 4.395 1.950 4.565 2.120 ;
        RECT 5.345 1.950 5.515 2.120 ;
        RECT 3.940 1.580 4.110 1.750 ;
        RECT 4.850 1.580 5.020 1.750 ;
        RECT 6.345 1.950 6.515 2.120 ;
        RECT 5.845 1.580 6.015 1.750 ;
        RECT 7.345 1.950 7.515 2.120 ;
        RECT 6.840 1.580 7.010 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__inv_16

#--------EOF---------

MACRO sky130_fd_sc_hs__maj3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__maj3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.570 3.715 0.670 ;
        RECT 2.645 0.255 3.715 0.570 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.430 1.685 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.285 1.760 2.755 1.780 ;
        RECT 2.285 1.430 3.575 1.760 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.485 1.370 3.775 1.450 ;
        RECT 0.040 1.290 3.810 1.370 ;
        RECT 0.005 0.245 3.810 1.290 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.538500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.850 0.490 2.980 ;
        RECT 0.085 1.180 0.255 1.850 ;
        RECT 0.085 0.480 0.445 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.660 1.950 0.990 3.245 ;
        RECT 1.565 2.120 1.895 2.940 ;
        RECT 2.435 2.290 2.840 3.245 ;
        RECT 3.395 2.120 3.725 2.940 ;
        RECT 1.565 1.950 3.725 2.120 ;
        RECT 0.425 1.350 0.785 1.680 ;
        RECT 0.615 1.260 0.785 1.350 ;
        RECT 1.895 1.260 2.065 1.950 ;
        RECT 3.395 1.930 3.725 1.950 ;
        RECT 0.615 1.090 3.700 1.260 ;
        RECT 0.615 0.085 0.990 0.910 ;
        RECT 1.480 0.580 1.810 1.090 ;
        RECT 2.305 0.740 2.850 0.910 ;
        RECT 3.370 0.840 3.700 1.090 ;
        RECT 2.305 0.085 2.475 0.740 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__maj3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__maj3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__maj3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.180 1.795 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 2.305 1.245 2.975 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 3.215 1.630 3.715 1.780 ;
        RECT 3.215 1.300 4.535 1.630 ;
        RECT 3.215 1.245 3.715 1.300 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 4.770 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
        RECT 1.875 1.555 3.825 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.820 0.915 2.980 ;
        RECT 0.555 1.130 0.725 1.820 ;
        RECT 0.555 0.350 0.895 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.135 1.820 0.385 3.245 ;
        RECT 1.085 2.120 1.780 3.245 ;
        RECT 1.965 2.120 2.785 2.755 ;
        RECT 3.485 2.290 3.815 3.245 ;
        RECT 4.355 2.120 4.685 2.860 ;
        RECT 1.965 1.950 4.685 2.120 ;
        RECT 1.085 1.780 2.135 1.950 ;
        RECT 4.355 1.820 4.685 1.950 ;
        RECT 1.085 1.650 1.255 1.780 ;
        RECT 0.895 1.320 1.255 1.650 ;
        RECT 0.135 0.085 0.385 1.130 ;
        RECT 1.965 1.075 2.135 1.780 ;
        RECT 4.330 1.075 4.660 1.130 ;
        RECT 1.075 0.085 1.795 1.010 ;
        RECT 1.965 0.905 4.660 1.075 ;
        RECT 1.965 0.350 2.760 0.905 ;
        RECT 3.340 0.085 3.840 0.680 ;
        RECT 4.330 0.350 4.660 0.905 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__maj3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__maj3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__maj3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 2.105 1.875 4.570 2.045 ;
        RECT 2.105 1.800 2.275 1.875 ;
        RECT 1.800 1.470 2.275 1.800 ;
        RECT 4.240 1.470 4.570 1.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.300 1.465 1.705 ;
        RECT 2.525 1.300 3.235 1.705 ;
        RECT 1.135 1.130 3.235 1.300 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.300 4.010 1.705 ;
        RECT 4.755 1.470 5.220 1.800 ;
        RECT 4.755 1.300 4.925 1.470 ;
        RECT 3.485 1.130 4.925 1.300 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.365 3.820 1.395 ;
        RECT 0.005 0.945 8.120 1.365 ;
        RECT 0.005 0.245 8.155 0.945 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 2.015 6.695 2.980 ;
        RECT 7.345 2.015 7.515 2.980 ;
        RECT 6.365 1.845 7.515 2.015 ;
        RECT 7.345 1.650 7.515 1.845 ;
        RECT 7.345 1.480 8.035 1.650 ;
        RECT 7.805 1.175 8.035 1.480 ;
        RECT 6.425 1.005 8.035 1.175 ;
        RECT 6.425 0.475 6.675 1.005 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.130 1.940 0.380 3.245 ;
        RECT 0.580 2.905 1.860 3.075 ;
        RECT 0.580 2.215 0.910 2.905 ;
        RECT 1.095 2.385 1.350 2.735 ;
        RECT 1.530 2.555 1.860 2.905 ;
        RECT 2.060 2.555 2.320 3.245 ;
        RECT 2.490 2.905 3.820 3.075 ;
        RECT 2.490 2.555 2.820 2.905 ;
        RECT 2.990 2.385 3.320 2.735 ;
        RECT 3.490 2.555 3.820 2.905 ;
        RECT 3.990 2.555 4.320 3.245 ;
        RECT 4.510 2.725 4.840 2.980 ;
        RECT 5.410 2.725 5.740 2.980 ;
        RECT 4.510 2.555 5.740 2.725 ;
        RECT 1.095 2.215 5.290 2.385 ;
        RECT 1.095 2.045 1.410 2.215 ;
        RECT 0.795 1.875 1.410 2.045 ;
        RECT 4.960 2.140 5.290 2.215 ;
        RECT 4.960 1.970 5.560 2.140 ;
        RECT 0.115 0.085 0.445 1.285 ;
        RECT 0.795 0.960 0.965 1.875 ;
        RECT 5.390 1.675 5.560 1.970 ;
        RECT 5.940 1.940 6.190 3.245 ;
        RECT 6.895 2.185 7.145 3.245 ;
        RECT 7.715 1.820 8.045 3.245 ;
        RECT 5.390 1.345 7.150 1.675 ;
        RECT 5.390 1.300 5.560 1.345 ;
        RECT 5.095 1.130 5.560 1.300 ;
        RECT 5.095 0.960 5.265 1.130 ;
        RECT 0.795 0.790 1.465 0.960 ;
        RECT 0.625 0.435 0.955 0.620 ;
        RECT 1.135 0.605 1.465 0.790 ;
        RECT 1.635 0.435 1.965 0.960 ;
        RECT 0.625 0.265 1.965 0.435 ;
        RECT 2.145 0.085 2.315 0.960 ;
        RECT 2.495 0.435 2.885 0.935 ;
        RECT 3.065 0.790 5.265 0.960 ;
        RECT 3.065 0.605 3.315 0.790 ;
        RECT 3.495 0.435 3.825 0.620 ;
        RECT 2.495 0.265 3.825 0.435 ;
        RECT 4.005 0.085 4.335 0.620 ;
        RECT 4.505 0.425 4.835 0.620 ;
        RECT 5.095 0.595 5.265 0.790 ;
        RECT 5.445 0.425 5.775 0.960 ;
        RECT 4.505 0.255 5.775 0.425 ;
        RECT 5.955 0.085 6.205 1.175 ;
        RECT 6.855 0.085 7.185 0.835 ;
        RECT 7.715 0.085 8.045 0.835 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__maj3_4

#--------EOF---------

MACRO sky130_fd_sc_hs__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.180 2.275 1.550 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.345 1.220 1.685 1.550 ;
        RECT 1.515 0.980 1.685 1.220 ;
        RECT 2.455 0.980 2.785 1.550 ;
        RECT 1.515 0.810 2.785 0.980 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.350 0.835 1.780 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.305 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.795 1.820 4.235 2.980 ;
        RECT 4.065 1.130 4.235 1.820 ;
        RECT 3.865 0.350 4.235 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.230 0.445 2.700 ;
        RECT 0.650 2.400 0.980 3.245 ;
        RECT 1.150 2.905 3.125 3.075 ;
        RECT 1.150 2.230 1.320 2.905 ;
        RECT 0.115 2.060 1.320 2.230 ;
        RECT 0.115 1.950 0.445 2.060 ;
        RECT 0.115 1.130 0.285 1.950 ;
        RECT 2.065 1.890 2.395 2.735 ;
        RECT 1.005 1.720 2.395 1.890 ;
        RECT 0.115 0.540 0.445 1.130 ;
        RECT 0.625 0.680 0.835 1.130 ;
        RECT 1.005 1.020 1.175 1.720 ;
        RECT 2.955 1.650 3.125 2.905 ;
        RECT 3.295 1.820 3.625 3.245 ;
        RECT 2.955 1.320 3.355 1.650 ;
        RECT 3.525 1.300 3.895 1.630 ;
        RECT 3.525 1.150 3.695 1.300 ;
        RECT 1.005 0.850 1.345 1.020 ;
        RECT 0.625 0.085 1.005 0.680 ;
        RECT 1.175 0.640 1.345 0.850 ;
        RECT 2.955 0.980 3.695 1.150 ;
        RECT 2.955 0.640 3.125 0.980 ;
        RECT 1.175 0.390 3.125 0.640 ;
        RECT 3.295 0.085 3.625 0.810 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__mux2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__mux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.180 1.195 1.550 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.450 2.385 1.780 ;
        RECT 2.215 1.300 2.385 1.450 ;
        RECT 3.125 1.300 3.455 1.460 ;
        RECT 2.215 1.130 3.455 1.300 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 1.050 2.870 1.240 ;
        RECT 3.830 1.050 5.275 1.240 ;
        RECT 0.060 0.245 5.275 1.050 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.965 0.770 4.665 2.140 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.115 2.905 1.905 3.075 ;
        RECT 0.115 1.825 0.445 2.905 ;
        RECT 0.620 2.140 0.840 2.725 ;
        RECT 1.015 2.480 1.345 2.735 ;
        RECT 1.575 2.650 1.905 2.905 ;
        RECT 2.075 2.650 2.405 3.245 ;
        RECT 2.575 2.480 2.825 2.980 ;
        RECT 3.870 2.650 4.210 3.245 ;
        RECT 4.780 2.650 5.165 3.245 ;
        RECT 1.015 2.310 2.825 2.480 ;
        RECT 2.995 2.310 5.165 2.480 ;
        RECT 2.995 2.140 3.165 2.310 ;
        RECT 0.620 1.970 3.165 2.140 ;
        RECT 0.620 1.820 1.535 1.970 ;
        RECT 1.365 1.010 1.535 1.820 ;
        RECT 3.335 1.800 3.795 2.140 ;
        RECT 2.555 1.630 3.795 1.800 ;
        RECT 2.555 1.470 2.885 1.630 ;
        RECT 0.170 0.460 0.500 1.010 ;
        RECT 0.670 0.680 1.535 1.010 ;
        RECT 1.715 0.960 2.045 1.130 ;
        RECT 1.715 0.790 3.170 0.960 ;
        RECT 3.625 0.940 3.795 1.630 ;
        RECT 4.835 1.300 5.165 2.310 ;
        RECT 2.420 0.460 2.750 0.620 ;
        RECT 0.170 0.290 2.750 0.460 ;
        RECT 3.000 0.085 3.170 0.790 ;
        RECT 3.340 0.770 3.795 0.940 ;
        RECT 3.340 0.350 3.670 0.770 ;
        RECT 3.840 0.085 4.230 0.600 ;
        RECT 4.835 0.085 5.165 1.130 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__mux2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.640 1.450 7.075 1.780 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 7.325 1.450 8.175 1.780 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.738000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 2.220 3.165 2.325 ;
        RECT 0.665 2.155 3.165 2.220 ;
        RECT 0.665 2.050 1.675 2.155 ;
        RECT 0.665 1.780 0.835 2.050 ;
        RECT 0.425 1.350 0.835 1.780 ;
        RECT 2.995 1.765 3.165 2.155 ;
        RECT 2.995 1.435 3.745 1.765 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.815 1.260 5.685 1.365 ;
        RECT 0.160 1.140 5.685 1.260 ;
        RECT 0.160 0.245 8.635 1.140 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
        RECT 0.850 1.575 2.930 1.660 ;
        RECT 0.850 1.470 1.690 1.575 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.576550 ;
    PORT
      LAYER li1 ;
        RECT 2.440 1.880 2.770 1.985 ;
        RECT 1.085 1.710 2.770 1.880 ;
        RECT 1.085 1.370 2.755 1.710 ;
        RECT 1.310 0.370 1.640 1.370 ;
        RECT 2.330 0.370 2.755 1.370 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.085 2.560 0.445 2.860 ;
        RECT 0.650 2.730 0.995 3.245 ;
        RECT 1.820 2.835 2.150 3.245 ;
        RECT 3.060 2.835 3.390 3.245 ;
        RECT 1.165 2.560 3.505 2.665 ;
        RECT 0.085 2.495 3.505 2.560 ;
        RECT 0.085 2.390 1.335 2.495 ;
        RECT 0.085 1.950 0.445 2.390 ;
        RECT 3.335 2.105 3.505 2.495 ;
        RECT 3.675 2.605 3.925 2.975 ;
        RECT 4.130 2.775 4.460 3.245 ;
        RECT 5.200 2.775 5.450 3.245 ;
        RECT 5.620 2.710 7.115 2.980 ;
        RECT 5.620 2.605 5.790 2.710 ;
        RECT 3.675 2.435 5.790 2.605 ;
        RECT 7.695 2.540 8.025 2.980 ;
        RECT 3.675 2.275 3.925 2.435 ;
        RECT 5.960 2.370 8.025 2.540 ;
        RECT 5.960 2.265 6.130 2.370 ;
        RECT 0.085 1.150 0.255 1.950 ;
        RECT 3.335 1.935 4.085 2.105 ;
        RECT 4.665 2.095 6.130 2.265 ;
        RECT 8.195 2.200 8.525 2.980 ;
        RECT 4.665 1.935 5.140 2.095 ;
        RECT 6.300 1.950 8.525 2.200 ;
        RECT 3.915 1.765 4.085 1.935 ;
        RECT 6.300 1.780 6.470 1.950 ;
        RECT 3.915 1.435 4.985 1.765 ;
        RECT 5.385 1.450 6.470 1.780 ;
        RECT 5.155 1.265 8.020 1.280 ;
        RECT 0.085 0.470 0.600 1.150 ;
        RECT 0.770 0.085 1.100 1.150 ;
        RECT 1.810 0.085 2.140 1.070 ;
        RECT 2.925 0.085 3.255 1.255 ;
        RECT 3.520 1.110 8.020 1.265 ;
        RECT 3.520 1.095 5.325 1.110 ;
        RECT 3.520 0.575 3.850 1.095 ;
        RECT 5.495 0.925 7.090 0.940 ;
        RECT 4.020 0.085 4.490 0.905 ;
        RECT 4.660 0.770 7.090 0.925 ;
        RECT 4.660 0.755 5.665 0.770 ;
        RECT 4.660 0.575 4.990 0.755 ;
        RECT 5.170 0.085 5.575 0.585 ;
        RECT 5.835 0.425 6.590 0.600 ;
        RECT 6.760 0.595 7.090 0.770 ;
        RECT 7.260 0.425 7.590 0.940 ;
        RECT 7.770 0.595 8.020 1.110 ;
        RECT 8.355 1.030 8.525 1.950 ;
        RECT 8.190 0.425 8.525 1.030 ;
        RECT 5.835 0.255 8.525 0.425 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__mux2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux2i_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 2.865 1.780 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.180 3.725 1.550 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.487500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.550 1.855 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.050 3.790 1.240 ;
        RECT 0.005 0.245 3.790 1.050 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.857700 ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.035 3.225 2.735 ;
        RECT 2.495 0.705 3.225 1.035 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.105 2.100 0.355 3.245 ;
        RECT 0.555 2.100 0.890 2.980 ;
        RECT 0.720 1.520 0.890 2.100 ;
        RECT 1.080 2.120 1.330 2.980 ;
        RECT 1.530 2.290 1.860 3.245 ;
        RECT 2.060 2.905 3.735 3.075 ;
        RECT 2.060 2.290 2.310 2.905 ;
        RECT 2.505 2.120 2.835 2.735 ;
        RECT 1.080 1.950 2.835 2.120 ;
        RECT 1.080 1.820 1.330 1.950 ;
        RECT 3.405 1.820 3.735 2.905 ;
        RECT 1.800 1.520 2.130 1.680 ;
        RECT 0.720 1.350 2.130 1.520 ;
        RECT 0.720 0.905 0.890 1.350 ;
        RECT 0.115 0.085 0.365 0.905 ;
        RECT 0.545 0.405 0.890 0.905 ;
        RECT 1.105 1.010 2.275 1.180 ;
        RECT 1.105 0.350 1.435 1.010 ;
        RECT 1.605 0.085 1.935 0.840 ;
        RECT 2.105 0.520 2.275 1.010 ;
        RECT 3.395 0.520 3.680 1.010 ;
        RECT 2.105 0.350 3.680 0.520 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__mux2i_1

#--------EOF---------

MACRO sky130_fd_sc_hs__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux2i_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.180 1.315 1.550 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.430 3.235 1.775 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.804000 ;
    PORT
      LAYER li1 ;
        RECT 4.350 1.840 5.810 2.010 ;
        RECT 3.485 1.430 4.675 1.840 ;
        RECT 5.480 1.350 5.810 1.840 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.630 1.240 2.180 1.295 ;
        RECT 3.030 1.240 6.235 1.360 ;
        RECT 0.010 0.245 6.235 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.040950 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.115 0.445 2.980 ;
        RECT 0.085 1.945 2.845 2.115 ;
        RECT 0.085 1.820 0.445 1.945 ;
        RECT 0.085 1.010 0.255 1.820 ;
        RECT 0.085 0.425 0.450 1.010 ;
        RECT 2.580 0.425 2.910 0.580 ;
        RECT 0.085 0.255 2.910 0.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.615 2.455 0.945 2.980 ;
        RECT 3.075 2.965 3.470 3.245 ;
        RECT 1.685 2.795 2.395 2.955 ;
        RECT 4.210 2.850 4.555 3.245 ;
        RECT 1.685 2.680 3.525 2.795 ;
        RECT 4.760 2.680 5.090 2.980 ;
        RECT 1.685 2.625 5.090 2.680 ;
        RECT 3.355 2.510 5.090 2.625 ;
        RECT 0.615 2.340 3.185 2.455 ;
        RECT 0.615 2.285 4.005 2.340 ;
        RECT 3.015 2.010 4.005 2.285 ;
        RECT 4.760 2.180 5.090 2.510 ;
        RECT 5.260 2.180 5.590 3.245 ;
        RECT 5.795 2.180 6.150 2.860 ;
        RECT 1.740 1.090 4.030 1.260 ;
        RECT 0.640 0.765 0.970 1.010 ;
        RECT 1.740 0.935 2.070 1.090 ;
        RECT 3.650 1.000 4.030 1.090 ;
        RECT 4.910 1.180 5.240 1.670 ;
        RECT 5.980 1.180 6.150 2.180 ;
        RECT 4.910 1.010 6.150 1.180 ;
        RECT 2.240 0.830 3.250 0.920 ;
        RECT 2.240 0.765 5.115 0.830 ;
        RECT 0.640 0.750 5.115 0.765 ;
        RECT 0.640 0.595 2.410 0.750 ;
        RECT 3.080 0.660 5.115 0.750 ;
        RECT 4.735 0.500 5.115 0.660 ;
        RECT 3.140 0.085 3.470 0.490 ;
        RECT 4.210 0.085 4.555 0.490 ;
        RECT 5.285 0.085 5.615 0.840 ;
        RECT 5.795 0.570 6.150 1.010 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__mux2i_2

#--------EOF---------

MACRO sky130_fd_sc_hs__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux2i_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.680 3.235 1.780 ;
        RECT 2.225 1.350 3.235 1.680 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.350 1.885 1.780 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.479000 ;
    PORT
      LAYER li1 ;
        RECT 7.080 1.180 9.475 1.540 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.745 1.295 6.200 1.360 ;
        RECT 0.005 1.280 6.200 1.295 ;
        RECT 0.005 0.245 9.935 1.280 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.868700 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.120 0.365 2.980 ;
        RECT 1.095 2.120 1.265 2.735 ;
        RECT 1.915 2.120 2.245 2.735 ;
        RECT 2.915 2.120 3.245 2.395 ;
        RECT 3.915 2.120 4.245 2.395 ;
        RECT 0.115 1.950 4.245 2.120 ;
        RECT 0.115 1.820 0.365 1.950 ;
        RECT 3.485 1.550 4.245 1.950 ;
        RECT 0.115 1.180 0.365 1.185 ;
        RECT 3.915 1.180 4.085 1.550 ;
        RECT 0.115 1.010 4.085 1.180 ;
        RECT 0.115 0.405 0.365 1.010 ;
        RECT 1.055 0.595 1.225 1.010 ;
        RECT 1.920 0.935 4.085 1.010 ;
        RECT 1.920 0.595 2.250 0.935 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.565 2.905 6.560 3.075 ;
        RECT 0.565 2.290 0.895 2.905 ;
        RECT 1.465 2.290 1.715 2.905 ;
        RECT 2.415 2.565 5.130 2.735 ;
        RECT 5.300 2.730 6.560 2.905 ;
        RECT 6.730 2.730 7.060 3.245 ;
        RECT 2.415 2.290 2.745 2.565 ;
        RECT 3.415 2.290 3.745 2.565 ;
        RECT 4.960 2.560 5.130 2.565 ;
        RECT 7.230 2.560 7.560 2.980 ;
        RECT 7.730 2.730 8.060 3.245 ;
        RECT 8.230 2.560 8.560 2.980 ;
        RECT 4.960 2.390 8.560 2.560 ;
        RECT 8.760 2.220 9.010 3.245 ;
        RECT 4.475 2.050 9.010 2.220 ;
        RECT 4.475 1.840 6.080 2.050 ;
        RECT 9.185 1.880 9.455 2.700 ;
        RECT 9.635 2.050 9.965 3.245 ;
        RECT 6.670 1.710 9.825 1.880 ;
        RECT 6.670 1.670 6.840 1.710 ;
        RECT 5.150 1.340 6.840 1.670 ;
        RECT 4.255 1.000 6.715 1.170 ;
        RECT 9.655 1.010 9.825 1.710 ;
        RECT 0.545 0.425 0.875 0.840 ;
        RECT 1.405 0.425 1.735 0.840 ;
        RECT 4.255 0.765 4.425 1.000 ;
        RECT 6.385 0.920 6.715 1.000 ;
        RECT 7.405 0.840 8.825 1.010 ;
        RECT 2.420 0.595 4.425 0.765 ;
        RECT 4.595 0.750 5.525 0.830 ;
        RECT 7.405 0.750 7.735 0.840 ;
        RECT 4.595 0.660 7.735 0.750 ;
        RECT 4.595 0.425 4.765 0.660 ;
        RECT 5.355 0.580 7.735 0.660 ;
        RECT 0.545 0.255 4.765 0.425 ;
        RECT 4.935 0.085 5.185 0.490 ;
        RECT 5.875 0.085 6.205 0.410 ;
        RECT 6.895 0.085 7.225 0.410 ;
        RECT 7.405 0.390 7.735 0.580 ;
        RECT 7.905 0.085 8.325 0.640 ;
        RECT 8.495 0.390 8.825 0.840 ;
        RECT 8.995 0.085 9.325 1.010 ;
        RECT 9.495 0.390 9.825 1.010 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__mux2i_4

#--------EOF---------

MACRO sky130_fd_sc_hs__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.990 1.215 1.320 1.780 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.000 1.215 3.330 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.500 1.215 3.870 2.150 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 5.850 1.445 6.180 1.780 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.738000 ;
    PORT
      LAYER li1 ;
        RECT 0.450 1.215 0.820 1.780 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 8.205 1.350 8.535 1.780 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.160 1.290 7.545 1.395 ;
        RECT 6.160 1.140 9.520 1.290 ;
        RECT 0.005 0.245 9.520 1.140 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
        RECT 0.680 1.525 4.260 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.558100 ;
    PORT
      LAYER li1 ;
        RECT 9.220 2.560 9.485 2.890 ;
        RECT 9.245 1.180 9.485 2.560 ;
        RECT 9.080 0.400 9.485 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.110 1.950 0.555 2.880 ;
        RECT 0.725 1.950 1.055 3.245 ;
        RECT 2.030 2.505 2.550 2.725 ;
        RECT 3.265 2.675 3.595 3.245 ;
        RECT 3.795 2.905 5.550 3.075 ;
        RECT 3.795 2.505 4.020 2.905 ;
        RECT 2.030 2.335 4.020 2.505 ;
        RECT 0.110 1.030 0.280 1.950 ;
        RECT 2.030 1.685 2.550 2.335 ;
        RECT 4.305 2.165 5.165 2.735 ;
        RECT 5.350 2.505 5.550 2.905 ;
        RECT 5.730 2.675 6.060 3.245 ;
        RECT 6.290 2.505 6.620 2.980 ;
        RECT 5.350 2.335 6.620 2.505 ;
        RECT 4.305 1.995 5.680 2.165 ;
        RECT 1.530 1.200 1.860 1.530 ;
        RECT 1.530 1.030 1.700 1.200 ;
        RECT 2.030 1.030 2.200 1.685 ;
        RECT 0.110 0.860 1.700 1.030 ;
        RECT 0.110 0.350 0.445 0.860 ;
        RECT 0.700 0.085 1.090 0.680 ;
        RECT 1.530 0.425 1.700 0.860 ;
        RECT 1.875 0.595 2.200 1.030 ;
        RECT 2.460 1.045 2.790 1.450 ;
        RECT 4.080 1.045 4.410 1.450 ;
        RECT 4.580 1.445 5.340 1.775 ;
        RECT 4.580 1.045 4.750 1.445 ;
        RECT 5.510 1.275 5.680 1.995 ;
        RECT 6.290 1.950 6.620 2.335 ;
        RECT 6.790 2.905 8.520 3.075 ;
        RECT 2.460 0.875 4.750 1.045 ;
        RECT 4.920 1.105 6.235 1.275 ;
        RECT 2.460 0.425 2.630 0.875 ;
        RECT 4.920 0.705 5.090 1.105 ;
        RECT 1.530 0.255 2.630 0.425 ;
        RECT 3.125 0.085 3.715 0.680 ;
        RECT 4.210 0.375 5.090 0.705 ;
        RECT 5.260 0.085 5.590 0.935 ;
        RECT 5.985 0.445 6.235 1.105 ;
        RECT 6.405 0.785 6.575 1.950 ;
        RECT 6.790 1.285 7.120 2.905 ;
        RECT 6.745 1.115 7.120 1.285 ;
        RECT 7.290 1.945 7.620 2.735 ;
        RECT 7.850 1.950 8.180 2.735 ;
        RECT 8.350 2.120 8.520 2.905 ;
        RECT 8.690 2.290 9.020 3.245 ;
        RECT 8.350 1.950 8.915 2.120 ;
        RECT 7.290 1.275 7.460 1.945 ;
        RECT 7.850 1.775 8.035 1.950 ;
        RECT 7.630 1.445 8.035 1.775 ;
        RECT 6.745 0.955 6.925 1.115 ;
        RECT 7.290 1.105 7.695 1.275 ;
        RECT 7.105 0.785 7.355 0.935 ;
        RECT 6.405 0.615 7.355 0.785 ;
        RECT 7.105 0.605 7.355 0.615 ;
        RECT 5.985 0.435 6.485 0.445 ;
        RECT 7.525 0.435 7.695 1.105 ;
        RECT 7.865 1.180 8.035 1.445 ;
        RECT 8.745 1.680 8.915 1.950 ;
        RECT 8.745 1.350 9.075 1.680 ;
        RECT 7.865 0.500 8.410 1.180 ;
        RECT 5.985 0.265 7.695 0.435 ;
        RECT 8.580 0.085 8.910 1.180 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
  END
END sky130_fd_sc_hs__mux4_1

#--------EOF---------

MACRO sky130_fd_sc_hs__mux4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.450 3.685 1.780 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.450 1.315 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 5.915 1.180 6.345 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.450 4.195 1.780 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.768000 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.280 0.805 1.550 ;
        RECT 1.485 1.280 1.845 1.590 ;
        RECT 0.435 1.260 1.845 1.280 ;
        RECT 2.835 1.280 3.105 1.780 ;
        RECT 4.395 1.280 4.725 1.550 ;
        RECT 5.475 1.280 5.745 1.750 ;
        RECT 0.435 1.180 1.655 1.260 ;
        RECT 0.635 1.110 1.655 1.180 ;
        RECT 1.485 0.590 1.655 1.110 ;
        RECT 2.835 1.110 5.745 1.280 ;
        RECT 2.835 0.590 3.105 1.110 ;
        RECT 1.485 0.420 3.105 0.590 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.507000 ;
    PORT
      LAYER li1 ;
        RECT 6.900 1.450 7.555 1.780 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.560 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.120 1.375 8.065 1.470 ;
        RECT 7.120 1.370 8.640 1.375 ;
        RECT 7.120 1.240 10.520 1.370 ;
        RECT 0.025 0.245 10.520 1.240 ;
        RECT 0.000 0.000 10.560 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.760 10.750 3.520 ;
        RECT -0.190 1.660 6.910 1.760 ;
        RECT 8.275 1.660 10.750 1.760 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.560 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 9.650 1.820 10.000 2.980 ;
        RECT 9.650 0.440 9.980 1.820 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.560 3.415 ;
        RECT 0.255 2.150 0.585 2.980 ;
        RECT 0.095 1.920 0.585 2.150 ;
        RECT 0.755 1.950 1.085 3.245 ;
        RECT 0.095 1.010 0.265 1.920 ;
        RECT 2.045 1.450 2.325 2.150 ;
        RECT 2.495 2.120 3.445 2.980 ;
        RECT 3.615 2.290 3.945 3.245 ;
        RECT 5.055 2.660 5.945 2.910 ;
        RECT 6.165 2.710 6.495 3.245 ;
        RECT 7.200 2.905 9.130 3.075 ;
        RECT 7.200 2.710 7.530 2.905 ;
        RECT 5.775 2.540 5.945 2.660 ;
        RECT 7.810 2.565 8.790 2.735 ;
        RECT 7.810 2.540 7.980 2.565 ;
        RECT 4.115 2.320 5.605 2.490 ;
        RECT 5.775 2.370 7.980 2.540 ;
        RECT 4.115 2.120 4.285 2.320 ;
        RECT 5.435 2.200 5.605 2.320 ;
        RECT 2.495 1.950 4.285 2.120 ;
        RECT 2.495 1.090 2.665 1.950 ;
        RECT 4.925 1.460 5.265 2.150 ;
        RECT 5.435 1.960 7.080 2.200 ;
        RECT 6.560 1.950 7.080 1.960 ;
        RECT 7.650 1.950 7.980 2.370 ;
        RECT 6.560 1.280 6.730 1.950 ;
        RECT 8.200 1.780 8.450 2.395 ;
        RECT 7.725 1.450 8.450 1.780 ;
        RECT 6.560 1.110 7.955 1.280 ;
        RECT 0.095 0.500 0.465 1.010 ;
        RECT 0.820 0.085 1.150 0.940 ;
        RECT 1.850 0.760 2.665 1.090 ;
        RECT 3.445 0.085 3.925 0.940 ;
        RECT 4.530 0.770 8.015 0.940 ;
        RECT 8.185 0.935 8.450 1.450 ;
        RECT 4.530 0.350 5.105 0.770 ;
        RECT 6.140 0.085 6.470 0.600 ;
        RECT 6.690 0.350 6.940 0.770 ;
        RECT 7.845 0.765 8.015 0.770 ;
        RECT 8.620 0.765 8.790 2.565 ;
        RECT 7.120 0.425 7.450 0.600 ;
        RECT 7.845 0.595 8.790 0.765 ;
        RECT 8.960 1.680 9.130 2.905 ;
        RECT 9.300 1.850 9.470 3.245 ;
        RECT 10.200 1.820 10.450 3.245 ;
        RECT 8.960 1.350 9.385 1.680 ;
        RECT 8.960 0.425 9.130 1.350 ;
        RECT 7.120 0.255 9.130 0.425 ;
        RECT 9.300 0.085 9.470 1.180 ;
        RECT 10.160 0.085 10.410 1.260 ;
        RECT 0.000 -0.085 10.560 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 0.155 1.950 0.325 2.120 ;
        RECT 2.075 1.950 2.245 2.120 ;
        RECT 4.955 1.950 5.125 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
      LAYER met1 ;
        RECT 0.095 2.105 0.385 2.150 ;
        RECT 2.015 2.105 2.305 2.150 ;
        RECT 4.895 2.105 5.185 2.150 ;
        RECT 0.095 1.965 5.185 2.105 ;
        RECT 0.095 1.920 0.385 1.965 ;
        RECT 2.015 1.920 2.305 1.965 ;
        RECT 4.895 1.920 5.185 1.965 ;
  END
END sky130_fd_sc_hs__mux4_2

#--------EOF---------

MACRO sky130_fd_sc_hs__mux4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__mux4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.470 2.355 1.800 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.890 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.260 9.475 1.775 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 9.725 1.445 10.435 1.775 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.263000 ;
    PORT
      LAYER li1 ;
        RECT 7.295 1.435 8.515 1.775 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.771000 ;
    PORT
      LAYER li1 ;
        RECT 12.150 1.300 12.835 1.780 ;
        RECT 13.540 1.300 13.865 1.550 ;
        RECT 12.150 1.275 13.865 1.300 ;
        RECT 12.665 1.130 13.865 1.275 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 16.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.365 2.420 1.400 ;
        RECT 0.005 1.240 4.825 1.365 ;
        RECT 5.825 1.240 8.175 1.375 ;
        RECT 0.005 1.140 8.175 1.240 ;
        RECT 13.795 1.140 16.795 1.240 ;
        RECT 0.005 0.245 16.795 1.140 ;
        RECT 0.000 0.000 16.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 16.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 14.875 1.970 15.205 2.980 ;
        RECT 15.825 1.970 16.155 2.980 ;
        RECT 14.875 1.800 16.675 1.970 ;
        RECT 16.445 1.130 16.675 1.800 ;
        RECT 15.065 0.960 16.675 1.130 ;
        RECT 15.065 0.350 15.315 0.960 ;
        RECT 15.925 0.350 16.175 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 16.800 3.415 ;
        RECT 0.115 1.950 0.365 3.245 ;
        RECT 0.565 2.140 0.895 2.980 ;
        RECT 1.095 2.310 1.345 3.245 ;
        RECT 1.515 2.480 1.845 2.980 ;
        RECT 2.045 2.650 2.295 3.245 ;
        RECT 2.525 2.905 4.720 3.075 ;
        RECT 2.525 2.650 2.860 2.905 ;
        RECT 3.045 2.480 3.300 2.735 ;
        RECT 1.515 2.310 3.300 2.480 ;
        RECT 0.565 1.970 2.695 2.140 ;
        RECT 0.565 1.950 0.895 1.970 ;
        RECT 2.525 1.770 2.695 1.970 ;
        RECT 2.990 1.940 3.300 2.310 ;
        RECT 3.490 1.940 3.820 2.905 ;
        RECT 4.020 1.770 4.190 2.735 ;
        RECT 2.525 1.600 4.190 1.770 ;
        RECT 4.375 1.920 4.720 2.905 ;
        RECT 2.525 1.300 4.205 1.430 ;
        RECT 0.115 1.030 1.370 1.280 ;
        RECT 0.115 0.085 0.365 1.030 ;
        RECT 0.545 0.470 0.875 0.860 ;
        RECT 1.045 0.640 1.370 1.030 ;
        RECT 1.550 1.260 4.205 1.300 ;
        RECT 1.550 1.130 2.695 1.260 ;
        RECT 1.550 0.960 1.800 1.130 ;
        RECT 3.050 0.960 3.380 1.090 ;
        RECT 1.970 0.790 3.380 0.960 ;
        RECT 1.575 0.620 2.140 0.790 ;
        RECT 1.575 0.470 1.810 0.620 ;
        RECT 0.545 0.275 1.810 0.470 ;
        RECT 1.980 0.085 2.310 0.450 ;
        RECT 2.540 0.425 2.870 0.620 ;
        RECT 3.050 0.595 3.380 0.790 ;
        RECT 3.605 0.425 3.775 1.090 ;
        RECT 3.955 0.595 4.205 1.260 ;
        RECT 4.375 1.180 4.545 1.920 ;
        RECT 4.950 1.680 5.200 2.980 ;
        RECT 5.400 1.820 5.730 3.245 ;
        RECT 6.410 2.905 8.150 3.075 ;
        RECT 8.320 2.965 8.650 3.245 ;
        RECT 9.390 2.965 9.730 3.245 ;
        RECT 5.960 2.035 6.210 2.905 ;
        RECT 6.410 2.205 6.740 2.905 ;
        RECT 7.980 2.795 8.150 2.905 ;
        RECT 9.935 2.795 10.265 2.980 ;
        RECT 6.940 2.115 7.125 2.735 ;
        RECT 7.310 2.455 7.640 2.735 ;
        RECT 7.980 2.625 10.265 2.795 ;
        RECT 7.310 2.285 9.185 2.455 ;
        RECT 9.935 2.285 10.265 2.625 ;
        RECT 10.465 2.285 10.635 3.245 ;
        RECT 10.805 2.905 12.975 3.075 ;
        RECT 10.805 2.115 10.975 2.905 ;
        RECT 6.940 2.035 10.975 2.115 ;
        RECT 5.960 1.945 10.975 2.035 ;
        RECT 11.145 2.565 12.475 2.735 ;
        RECT 5.960 1.865 7.125 1.945 ;
        RECT 4.715 1.535 5.200 1.680 ;
        RECT 6.035 1.535 6.705 1.695 ;
        RECT 4.715 1.365 6.705 1.535 ;
        RECT 4.715 1.350 5.200 1.365 ;
        RECT 4.375 0.425 4.715 1.180 ;
        RECT 2.540 0.255 4.715 0.425 ;
        RECT 4.945 0.350 5.200 1.350 ;
        RECT 6.940 1.265 7.125 1.865 ;
        RECT 6.875 1.195 7.125 1.265 ;
        RECT 5.375 0.085 5.705 1.130 ;
        RECT 5.935 1.025 7.125 1.195 ;
        RECT 5.935 0.585 6.185 1.025 ;
        RECT 6.365 0.425 6.695 0.855 ;
        RECT 6.875 0.765 7.125 1.025 ;
        RECT 7.305 1.095 8.325 1.265 ;
        RECT 7.305 0.935 7.555 1.095 ;
        RECT 8.155 1.090 8.325 1.095 ;
        RECT 7.735 0.765 7.985 0.925 ;
        RECT 8.155 0.920 10.115 1.090 ;
        RECT 6.875 0.595 7.985 0.765 ;
        RECT 8.155 0.580 9.255 0.750 ;
        RECT 8.155 0.425 8.325 0.580 ;
        RECT 6.365 0.255 8.325 0.425 ;
        RECT 8.495 0.085 8.825 0.410 ;
        RECT 9.005 0.350 9.255 0.580 ;
        RECT 9.435 0.085 9.685 0.750 ;
        RECT 9.865 0.350 10.115 0.920 ;
        RECT 10.295 0.085 10.545 1.030 ;
        RECT 10.715 0.425 10.885 1.945 ;
        RECT 11.145 1.030 11.475 2.565 ;
        RECT 11.055 0.765 11.475 1.030 ;
        RECT 11.645 1.105 11.975 2.395 ;
        RECT 12.145 2.230 12.475 2.565 ;
        RECT 12.645 2.400 12.975 2.905 ;
        RECT 13.145 2.230 13.475 2.980 ;
        RECT 12.145 2.060 13.475 2.230 ;
        RECT 12.145 1.950 12.475 2.060 ;
        RECT 13.875 1.890 14.205 2.980 ;
        RECT 13.005 1.720 14.205 1.890 ;
        RECT 14.375 1.820 14.705 3.245 ;
        RECT 15.405 2.140 15.655 3.245 ;
        RECT 16.325 2.140 16.655 3.245 ;
        RECT 13.005 1.470 13.330 1.720 ;
        RECT 11.645 0.960 12.495 1.105 ;
        RECT 14.035 0.960 14.205 1.720 ;
        RECT 11.645 0.935 13.175 0.960 ;
        RECT 12.325 0.790 13.175 0.935 ;
        RECT 11.055 0.620 12.155 0.765 ;
        RECT 11.055 0.595 12.675 0.620 ;
        RECT 12.860 0.595 13.175 0.790 ;
        RECT 11.985 0.425 12.675 0.595 ;
        RECT 13.345 0.425 13.675 0.960 ;
        RECT 13.905 0.595 14.205 0.960 ;
        RECT 14.375 1.300 16.210 1.630 ;
        RECT 14.375 0.425 14.545 1.300 ;
        RECT 10.715 0.255 11.815 0.425 ;
        RECT 11.985 0.255 14.545 0.425 ;
        RECT 14.715 0.085 14.885 1.130 ;
        RECT 15.495 0.085 15.745 0.790 ;
        RECT 16.355 0.085 16.685 0.790 ;
        RECT 0.000 -0.085 16.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 4.475 1.950 4.645 2.120 ;
        RECT 11.675 1.950 11.845 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
      LAYER met1 ;
        RECT 4.415 2.105 4.705 2.150 ;
        RECT 11.615 2.105 11.905 2.150 ;
        RECT 4.415 1.965 11.905 2.105 ;
        RECT 4.415 1.920 4.705 1.965 ;
        RECT 11.615 1.920 11.905 1.965 ;
  END
END sky130_fd_sc_hs__mux4_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.180 1.335 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 1.390 1.240 ;
        RECT 0.000 0.000 1.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.440 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.546900 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.180 0.835 2.980 ;
        RECT 0.665 1.010 0.835 1.180 ;
        RECT 0.665 0.840 1.280 1.010 ;
        RECT 0.950 0.350 1.280 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.440 3.415 ;
        RECT 0.105 1.820 0.435 3.245 ;
        RECT 1.005 1.820 1.335 3.245 ;
        RECT 0.130 0.085 0.460 1.010 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
  END
END sky130_fd_sc_hs__nand2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.350 1.815 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 1.315 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.916200 ;
    PORT
      LAYER li1 ;
        RECT 0.570 2.120 0.820 2.980 ;
        RECT 1.560 2.120 1.730 2.980 ;
        RECT 0.570 1.950 2.275 2.120 ;
        RECT 2.045 1.180 2.275 1.950 ;
        RECT 1.455 1.010 2.275 1.180 ;
        RECT 1.455 0.595 1.785 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.120 1.820 0.370 3.245 ;
        RECT 1.020 2.290 1.350 3.245 ;
        RECT 1.930 2.290 2.260 3.245 ;
        RECT 0.115 1.010 1.275 1.180 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.105 0.425 1.275 1.010 ;
        RECT 1.955 0.425 2.285 0.840 ;
        RECT 1.105 0.255 2.285 0.425 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__nand2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.350 3.795 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.680 2.275 1.780 ;
        RECT 0.510 1.350 2.275 1.680 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.286100 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 1.660 2.980 ;
        RECT 2.330 2.120 3.705 2.980 ;
        RECT 0.615 1.950 4.195 2.120 ;
        RECT 3.965 1.180 4.195 1.950 ;
        RECT 2.335 1.010 4.195 1.180 ;
        RECT 2.335 0.610 2.665 1.010 ;
        RECT 3.335 0.610 3.705 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 1.850 0.445 3.245 ;
        RECT 1.830 2.290 2.160 3.245 ;
        RECT 3.875 2.290 4.205 3.245 ;
        RECT 0.115 1.010 2.165 1.180 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.805 ;
        RECT 1.055 0.350 1.225 1.010 ;
        RECT 1.405 0.085 1.735 0.805 ;
        RECT 1.915 0.425 2.165 1.010 ;
        RECT 2.835 0.425 3.165 0.805 ;
        RECT 3.875 0.425 4.205 0.805 ;
        RECT 1.915 0.255 4.205 0.425 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__nand2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.550 7.555 1.780 ;
        RECT 5.185 1.220 7.555 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 4.195 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.790 8.110 1.240 ;
        RECT 0.005 0.245 8.155 0.790 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.284800 ;
    PORT
      LAYER li1 ;
        RECT 2.140 2.120 2.470 2.980 ;
        RECT 4.380 2.120 4.710 2.980 ;
        RECT 2.140 1.950 4.710 2.120 ;
        RECT 5.940 2.120 6.270 2.980 ;
        RECT 7.320 2.120 7.550 2.980 ;
        RECT 5.940 1.950 7.895 2.120 ;
        RECT 4.380 1.130 4.710 1.950 ;
        RECT 4.335 1.050 4.710 1.130 ;
        RECT 7.725 1.050 7.895 1.950 ;
        RECT 4.335 0.770 7.895 1.050 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.660 1.950 1.970 3.245 ;
        RECT 2.640 2.290 4.210 3.245 ;
        RECT 4.880 1.820 5.210 3.245 ;
        RECT 5.440 1.820 5.770 3.245 ;
        RECT 6.440 2.290 7.150 3.245 ;
        RECT 7.720 2.290 8.050 3.245 ;
        RECT 0.105 1.180 1.860 1.355 ;
        RECT 0.105 1.165 4.155 1.180 ;
        RECT 0.105 0.350 0.355 1.165 ;
        RECT 1.035 1.010 4.155 1.165 ;
        RECT 0.535 0.085 0.865 0.995 ;
        RECT 1.035 0.350 1.225 1.010 ;
        RECT 1.395 0.085 1.725 0.840 ;
        RECT 1.895 0.350 2.155 1.010 ;
        RECT 2.325 0.085 2.905 0.840 ;
        RECT 3.075 0.350 3.305 1.010 ;
        RECT 3.475 0.085 3.805 0.840 ;
        RECT 3.985 0.600 4.155 1.010 ;
        RECT 3.985 0.350 8.045 0.600 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__nand2_8

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.835 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.350 1.345 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.295 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.710200 ;
    PORT
      LAYER li1 ;
        RECT 1.085 2.460 1.565 2.980 ;
        RECT 1.085 2.290 2.255 2.460 ;
        RECT 2.085 1.130 2.255 2.290 ;
        RECT 1.855 0.350 2.255 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.115 2.120 0.445 2.700 ;
        RECT 0.650 2.290 0.915 3.245 ;
        RECT 1.735 2.650 2.070 3.245 ;
        RECT 0.115 1.950 1.685 2.120 ;
        RECT 1.515 1.630 1.685 1.950 ;
        RECT 1.515 1.300 1.915 1.630 ;
        RECT 1.515 1.130 1.685 1.300 ;
        RECT 0.115 0.960 1.685 1.130 ;
        RECT 0.115 0.540 0.380 0.960 ;
        RECT 0.550 0.085 1.220 0.790 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__nand2b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.570 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.350 2.775 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.115 1.140 3.355 1.240 ;
        RECT 0.005 0.245 3.355 1.140 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.879200 ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.950 2.795 2.200 ;
        RECT 1.645 1.820 2.275 1.950 ;
        RECT 2.045 1.390 2.275 1.820 ;
        RECT 1.700 1.220 2.275 1.390 ;
        RECT 1.700 0.630 1.870 1.220 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.120 0.445 2.860 ;
        RECT 0.725 2.290 1.095 3.245 ;
        RECT 2.015 2.710 2.345 3.245 ;
        RECT 2.915 2.710 3.245 3.245 ;
        RECT 1.305 2.370 3.245 2.540 ;
        RECT 0.115 1.950 0.975 2.120 ;
        RECT 0.805 1.470 0.975 1.950 ;
        RECT 0.805 1.180 1.135 1.470 ;
        RECT 0.115 1.140 1.135 1.180 ;
        RECT 0.115 1.010 0.975 1.140 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 1.305 0.970 1.475 2.370 ;
        RECT 3.075 1.130 3.245 2.370 ;
        RECT 0.615 0.085 0.875 0.840 ;
        RECT 1.190 0.425 1.520 0.970 ;
        RECT 2.050 0.425 2.380 1.050 ;
        RECT 1.190 0.255 2.380 0.425 ;
        RECT 2.560 0.085 2.730 1.130 ;
        RECT 2.915 0.350 3.245 1.130 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__nand2b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 1.115 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.630 5.655 1.780 ;
        RECT 3.845 1.300 5.655 1.630 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.634300 ;
    PORT
      LAYER li1 ;
        RECT 2.265 2.150 2.875 2.980 ;
        RECT 4.815 2.150 5.145 2.980 ;
        RECT 2.265 1.950 5.145 2.150 ;
        RECT 2.265 1.850 4.195 1.950 ;
        RECT 3.285 1.260 3.655 1.850 ;
        RECT 1.625 1.090 3.655 1.260 ;
        RECT 1.625 0.635 1.885 1.090 ;
        RECT 2.555 0.635 2.880 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.435 1.950 1.060 3.245 ;
        RECT 1.230 1.950 1.560 2.700 ;
        RECT 1.285 1.680 1.455 1.950 ;
        RECT 1.765 1.850 2.095 3.245 ;
        RECT 3.045 2.320 4.645 3.245 ;
        RECT 5.315 1.950 5.600 3.245 ;
        RECT 1.285 1.430 3.075 1.680 ;
        RECT 1.285 1.130 1.455 1.430 ;
        RECT 0.135 0.960 1.455 1.130 ;
        RECT 3.980 0.960 5.645 1.130 ;
        RECT 0.135 0.350 0.385 0.960 ;
        RECT 3.980 0.920 4.310 0.960 ;
        RECT 0.565 0.085 0.895 0.790 ;
        RECT 1.195 0.425 1.455 0.790 ;
        RECT 2.055 0.425 2.385 0.920 ;
        RECT 3.050 0.750 4.310 0.920 ;
        RECT 3.050 0.425 3.380 0.750 ;
        RECT 1.195 0.255 3.380 0.425 ;
        RECT 3.550 0.085 3.880 0.580 ;
        RECT 4.050 0.330 4.310 0.750 ;
        RECT 4.480 0.085 5.145 0.790 ;
        RECT 5.315 0.350 5.645 0.960 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__nand2b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.180 1.915 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.440 1.345 1.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.835 1.550 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 0.245 2.150 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.877300 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.890 1.045 2.980 ;
        RECT 1.735 1.890 2.255 2.980 ;
        RECT 0.605 1.720 2.255 1.890 ;
        RECT 2.085 1.010 2.255 1.720 ;
        RECT 1.710 0.840 2.255 1.010 ;
        RECT 1.710 0.350 2.040 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.185 1.820 0.435 3.245 ;
        RECT 1.215 2.060 1.545 3.245 ;
        RECT 0.320 0.085 0.650 1.010 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__nand3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.430 2.295 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.425 1.950 2.825 2.120 ;
        RECT 1.425 1.680 1.795 1.950 ;
        RECT 1.265 1.550 1.795 1.680 ;
        RECT 2.655 1.650 2.825 1.950 ;
        RECT 1.265 1.430 1.595 1.550 ;
        RECT 2.655 1.320 3.065 1.650 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.735 1.550 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.440 1.240 3.355 1.295 ;
        RECT 0.005 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.220800 ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.460 0.895 2.980 ;
        RECT 1.515 2.460 1.845 2.980 ;
        RECT 2.525 2.460 2.795 2.980 ;
        RECT 0.565 2.290 2.795 2.460 ;
        RECT 0.565 1.820 1.095 2.290 ;
        RECT 0.925 1.260 1.095 1.820 ;
        RECT 0.925 1.090 2.275 1.260 ;
        RECT 1.945 0.935 2.275 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.065 2.630 1.315 3.245 ;
        RECT 2.015 2.630 2.345 3.245 ;
        RECT 2.995 1.820 3.245 3.245 ;
        RECT 0.100 0.920 0.430 1.010 ;
        RECT 0.100 0.765 1.370 0.920 ;
        RECT 2.930 0.765 3.260 1.150 ;
        RECT 0.100 0.750 3.260 0.765 ;
        RECT 0.100 0.350 0.350 0.750 ;
        RECT 1.040 0.595 3.260 0.750 ;
        RECT 0.530 0.085 0.860 0.580 ;
        RECT 1.040 0.330 1.210 0.595 ;
        RECT 1.455 0.255 2.765 0.425 ;
        RECT 2.945 0.405 3.260 0.595 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__nand3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.350 1.535 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 2.560 1.630 3.715 1.780 ;
        RECT 2.130 1.350 3.715 1.630 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 4.495 1.630 6.115 1.780 ;
        RECT 4.140 1.340 6.115 1.630 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.950 6.235 1.280 ;
        RECT 0.005 0.245 6.235 0.950 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.004800 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 1.365 2.980 ;
        RECT 2.035 2.120 2.365 2.980 ;
        RECT 3.960 2.120 4.290 2.980 ;
        RECT 0.125 1.950 4.290 2.120 ;
        RECT 0.125 1.180 0.355 1.950 ;
        RECT 2.035 1.820 2.365 1.950 ;
        RECT 3.960 1.820 4.290 1.950 ;
        RECT 0.125 1.010 1.725 1.180 ;
        RECT 0.535 0.595 0.865 1.010 ;
        RECT 1.395 0.595 1.725 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.115 2.290 0.445 3.245 ;
        RECT 1.535 2.290 1.865 3.245 ;
        RECT 2.535 2.290 3.790 3.245 ;
        RECT 4.460 1.950 5.765 3.245 ;
        RECT 0.105 0.425 0.355 0.840 ;
        RECT 1.045 0.425 1.215 0.840 ;
        RECT 1.905 0.425 2.075 1.170 ;
        RECT 2.255 0.920 5.625 1.170 ;
        RECT 2.255 0.595 2.585 0.920 ;
        RECT 2.755 0.425 2.945 0.750 ;
        RECT 3.115 0.595 3.445 0.920 ;
        RECT 3.615 0.425 3.875 0.750 ;
        RECT 0.105 0.255 3.875 0.425 ;
        RECT 4.085 0.085 4.415 0.750 ;
        RECT 4.585 0.390 4.775 0.920 ;
        RECT 4.945 0.085 5.275 0.750 ;
        RECT 5.455 0.390 5.625 0.920 ;
        RECT 5.805 0.085 6.135 1.170 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__nand3_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.350 0.835 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 1.915 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.350 1.345 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.865 1.260 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006800 ;
    PORT
      LAYER li1 ;
        RECT 1.305 2.120 1.635 2.980 ;
        RECT 2.305 2.120 2.795 2.980 ;
        RECT 1.305 1.950 2.795 2.120 ;
        RECT 2.305 1.820 2.795 1.950 ;
        RECT 2.625 1.150 2.795 1.820 ;
        RECT 2.425 0.790 2.795 1.150 ;
        RECT 2.250 0.370 2.795 0.790 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.105 1.950 0.600 2.700 ;
        RECT 0.805 1.950 1.135 3.245 ;
        RECT 1.805 2.290 2.135 3.245 ;
        RECT 0.105 1.150 0.275 1.950 ;
        RECT 2.085 1.320 2.455 1.650 ;
        RECT 2.085 1.150 2.255 1.320 ;
        RECT 0.105 0.980 2.255 1.150 ;
        RECT 0.105 0.560 0.375 0.980 ;
        RECT 0.545 0.085 1.220 0.810 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__nand3b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.550 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 4.195 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.430 1.795 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.965 1.240 4.315 1.370 ;
        RECT 0.005 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.332800 ;
    PORT
      LAYER li1 ;
        RECT 1.260 2.120 1.635 2.980 ;
        RECT 2.335 2.120 2.585 2.980 ;
        RECT 3.365 2.120 3.695 2.980 ;
        RECT 1.260 1.950 3.695 2.120 ;
        RECT 2.525 1.180 2.800 1.950 ;
        RECT 2.470 1.010 2.800 1.180 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.305 2.120 0.635 2.980 ;
        RECT 0.830 2.290 1.075 3.245 ;
        RECT 1.805 2.290 2.135 3.245 ;
        RECT 2.790 2.290 3.120 3.245 ;
        RECT 0.305 1.950 0.890 2.120 ;
        RECT 3.875 1.950 4.205 3.245 ;
        RECT 0.720 1.260 0.890 1.950 ;
        RECT 2.025 1.350 2.355 1.680 ;
        RECT 2.025 1.260 2.195 1.350 ;
        RECT 0.100 1.090 2.195 1.260 ;
        RECT 0.100 0.450 0.350 1.090 ;
        RECT 0.530 0.085 0.820 0.910 ;
        RECT 1.005 0.840 2.105 0.920 ;
        RECT 2.970 0.840 3.790 1.180 ;
        RECT 1.005 0.750 3.790 0.840 ;
        RECT 1.005 0.330 1.255 0.750 ;
        RECT 1.935 0.670 3.790 0.750 ;
        RECT 1.435 0.085 1.765 0.580 ;
        RECT 3.960 0.500 4.220 1.180 ;
        RECT 1.975 0.330 4.220 0.500 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__nand3b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.350 1.095 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 5.820 1.180 7.075 1.650 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.350 3.235 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.315 1.240 3.545 1.280 ;
        RECT 0.315 0.860 7.640 1.240 ;
        RECT 0.315 0.245 7.675 0.860 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.866500 ;
    PORT
      LAYER li1 ;
        RECT 2.685 1.950 5.850 2.140 ;
        RECT 3.750 1.820 5.850 1.950 ;
        RECT 4.925 1.130 5.155 1.820 ;
        RECT 4.130 0.800 5.345 1.130 ;
        RECT 4.925 0.770 5.345 0.800 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.115 2.290 0.445 3.245 ;
        RECT 1.490 2.650 2.565 3.245 ;
        RECT 3.135 2.650 3.630 3.245 ;
        RECT 4.580 2.650 5.400 3.245 ;
        RECT 5.970 2.650 7.565 3.245 ;
        RECT 0.615 2.310 6.230 2.480 ;
        RECT 0.615 2.120 0.785 2.310 ;
        RECT 0.085 1.950 0.785 2.120 ;
        RECT 0.955 1.950 1.435 2.140 ;
        RECT 0.085 0.750 0.255 1.950 ;
        RECT 1.265 1.180 1.435 1.950 ;
        RECT 6.060 1.990 6.230 2.310 ;
        RECT 6.400 2.160 7.565 2.650 ;
        RECT 6.060 1.820 7.415 1.990 ;
        RECT 3.600 1.300 4.610 1.630 ;
        RECT 3.600 1.180 3.770 1.300 ;
        RECT 0.425 1.010 3.770 1.180 ;
        RECT 7.245 1.010 7.415 1.820 ;
        RECT 0.425 0.920 0.755 1.010 ;
        RECT 5.945 0.840 7.415 1.010 ;
        RECT 1.460 0.750 2.970 0.840 ;
        RECT 0.085 0.670 2.970 0.750 ;
        RECT 0.085 0.580 1.790 0.670 ;
        RECT 0.935 0.085 1.280 0.410 ;
        RECT 1.460 0.390 1.790 0.580 ;
        RECT 1.970 0.085 2.460 0.500 ;
        RECT 2.640 0.390 2.970 0.670 ;
        RECT 3.140 0.085 3.470 0.840 ;
        RECT 3.700 0.600 4.030 0.630 ;
        RECT 5.515 0.600 7.565 0.670 ;
        RECT 3.700 0.350 7.565 0.600 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__nand3b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.180 2.775 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.180 2.275 1.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.180 1.475 1.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.180 0.905 1.550 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.375 1.120 2.830 1.240 ;
        RECT 0.375 0.790 2.850 1.120 ;
        RECT 0.005 0.245 2.850 0.790 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.936500 ;
    PORT
      LAYER li1 ;
        RECT 0.875 2.150 1.205 2.980 ;
        RECT 1.935 2.150 2.265 2.980 ;
        RECT 0.875 1.890 2.265 2.150 ;
        RECT 0.235 1.820 2.265 1.890 ;
        RECT 0.235 1.720 1.205 1.820 ;
        RECT 0.235 1.010 0.405 1.720 ;
        RECT 0.235 0.840 2.740 1.010 ;
        RECT 2.410 0.350 2.740 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.375 2.060 0.705 3.245 ;
        RECT 1.400 2.320 1.730 3.245 ;
        RECT 2.435 1.820 2.765 3.245 ;
        RECT 0.110 0.085 0.785 0.600 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__nand4_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.350 4.215 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.680 1.350 3.715 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.430 1.350 2.440 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.090 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.950 4.700 1.240 ;
        RECT 0.005 0.245 4.785 0.950 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.633200 ;
    PORT
      LAYER li1 ;
        RECT 0.635 2.120 0.900 2.980 ;
        RECT 1.570 2.120 1.900 2.980 ;
        RECT 2.830 2.120 3.160 2.980 ;
        RECT 3.840 2.150 4.125 2.980 ;
        RECT 3.840 2.120 4.675 2.150 ;
        RECT 0.635 1.950 4.675 2.120 ;
        RECT 4.445 1.180 4.675 1.950 ;
        RECT 3.845 1.010 4.675 1.180 ;
        RECT 3.845 0.645 4.175 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 1.950 0.450 3.245 ;
        RECT 1.070 2.290 1.400 3.245 ;
        RECT 2.080 2.290 2.650 3.245 ;
        RECT 3.330 2.290 3.660 3.245 ;
        RECT 4.295 2.320 4.625 3.245 ;
        RECT 0.115 1.010 1.315 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.145 0.425 1.315 1.010 ;
        RECT 1.495 1.010 3.315 1.180 ;
        RECT 1.495 0.595 1.825 1.010 ;
        RECT 1.995 0.425 2.325 0.840 ;
        RECT 1.145 0.255 2.325 0.425 ;
        RECT 2.555 0.425 2.815 0.840 ;
        RECT 2.985 0.645 3.315 1.010 ;
        RECT 3.485 0.425 3.675 1.130 ;
        RECT 4.345 0.425 4.675 0.840 ;
        RECT 2.555 0.255 4.675 0.425 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__nand4_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 6.735 1.350 8.085 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 6.160 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 4.195 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 2.275 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.820 8.600 1.240 ;
        RECT 0.005 0.245 8.635 0.820 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.321600 ;
    PORT
      LAYER li1 ;
        RECT 1.820 2.120 2.150 2.980 ;
        RECT 2.820 2.120 3.430 2.980 ;
        RECT 4.670 2.120 5.280 2.980 ;
        RECT 7.320 2.120 8.010 2.980 ;
        RECT 1.820 1.950 8.515 2.120 ;
        RECT 8.285 1.130 8.515 1.950 ;
        RECT 6.745 0.880 8.515 1.130 ;
        RECT 6.815 0.800 7.005 0.880 ;
        RECT 7.755 0.800 7.945 0.880 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.115 1.950 1.650 3.245 ;
        RECT 2.320 2.290 2.650 3.245 ;
        RECT 3.600 2.290 4.500 3.245 ;
        RECT 5.450 2.290 7.140 3.245 ;
        RECT 8.190 2.290 8.520 3.245 ;
        RECT 0.115 1.010 2.575 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.115 0.350 1.445 1.010 ;
        RECT 1.615 0.085 1.945 0.840 ;
        RECT 2.245 0.680 2.575 1.010 ;
        RECT 2.745 0.880 6.215 1.130 ;
        RECT 2.745 0.850 3.935 0.880 ;
        RECT 5.095 0.800 5.285 0.880 ;
        RECT 5.955 0.800 6.145 0.880 ;
        RECT 2.245 0.350 4.365 0.680 ;
        RECT 4.595 0.520 4.925 0.710 ;
        RECT 5.455 0.520 5.785 0.710 ;
        RECT 6.315 0.520 6.645 0.710 ;
        RECT 7.175 0.520 7.505 0.710 ;
        RECT 8.195 0.520 8.525 0.710 ;
        RECT 4.595 0.350 8.525 0.520 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__nand4_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.180 0.815 1.550 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.395 1.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.180 1.855 1.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.180 1.315 1.550 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.345 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.012400 ;
    PORT
      LAYER li1 ;
        RECT 1.285 2.150 1.615 2.980 ;
        RECT 2.285 2.150 2.635 2.980 ;
        RECT 1.285 1.890 2.635 2.150 ;
        RECT 1.285 1.820 3.275 1.890 ;
        RECT 1.615 1.720 3.275 1.820 ;
        RECT 3.105 1.050 3.275 1.720 ;
        RECT 2.905 0.350 3.275 1.050 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.105 1.820 0.580 2.700 ;
        RECT 0.785 1.820 1.115 3.245 ;
        RECT 1.785 2.320 2.115 3.245 ;
        RECT 2.805 2.060 3.135 3.245 ;
        RECT 0.105 1.010 0.275 1.820 ;
        RECT 2.565 1.220 2.935 1.550 ;
        RECT 2.565 1.010 2.735 1.220 ;
        RECT 0.105 0.840 2.735 1.010 ;
        RECT 0.105 0.680 0.650 0.840 ;
        RECT 0.855 0.085 1.185 0.670 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__nand4b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.985 1.510 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.590 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.195 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 5.635 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.465 1.240 5.755 1.290 ;
        RECT 1.030 1.140 5.755 1.240 ;
        RECT 0.005 0.245 5.755 1.140 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.573400 ;
    PORT
      LAYER li1 ;
        RECT 1.550 2.120 1.825 2.980 ;
        RECT 2.760 2.120 3.090 2.980 ;
        RECT 3.760 2.120 4.090 2.980 ;
        RECT 4.860 2.120 5.190 2.980 ;
        RECT 1.550 1.950 5.190 2.120 ;
        RECT 1.550 1.850 1.825 1.950 ;
        RECT 2.760 1.820 3.235 1.950 ;
        RECT 3.005 1.180 3.235 1.820 ;
        RECT 1.535 1.010 3.235 1.180 ;
        RECT 1.535 0.800 1.895 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.505 1.850 0.835 2.860 ;
        RECT 1.040 2.020 1.370 3.245 ;
        RECT 1.995 2.290 2.590 3.245 ;
        RECT 3.260 2.290 3.590 3.245 ;
        RECT 4.320 2.290 4.650 3.245 ;
        RECT 5.360 1.950 5.645 3.245 ;
        RECT 0.505 1.680 1.325 1.850 ;
        RECT 1.155 1.350 1.720 1.680 ;
        RECT 1.155 1.010 1.325 1.350 ;
        RECT 0.115 0.840 1.325 1.010 ;
        RECT 3.575 0.930 5.645 1.180 ;
        RECT 0.115 0.350 0.365 0.840 ;
        RECT 2.075 0.670 3.345 0.840 ;
        RECT 0.545 0.085 0.875 0.670 ;
        RECT 2.075 0.630 2.325 0.670 ;
        RECT 1.105 0.350 2.325 0.630 ;
        RECT 3.015 0.595 3.345 0.670 ;
        RECT 3.575 0.595 3.825 0.930 ;
        RECT 2.505 0.425 2.835 0.500 ;
        RECT 4.005 0.425 4.335 0.760 ;
        RECT 2.505 0.255 4.335 0.425 ;
        RECT 4.505 0.400 4.695 0.930 ;
        RECT 4.865 0.085 5.195 0.760 ;
        RECT 5.395 0.400 5.645 0.930 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__nand4b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.835 1.780 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 3.130 1.430 4.140 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.350 7.555 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.300 9.015 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 9.115 1.240 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.665600 ;
    PORT
      LAYER li1 ;
        RECT 2.050 2.120 2.670 2.980 ;
        RECT 4.370 2.120 4.590 2.980 ;
        RECT 6.065 2.120 6.660 2.980 ;
        RECT 8.215 2.120 8.505 2.980 ;
        RECT 2.050 1.950 8.505 2.120 ;
        RECT 2.050 1.850 2.680 1.950 ;
        RECT 4.310 1.820 4.675 1.950 ;
        RECT 4.445 1.260 4.675 1.820 ;
        RECT 2.395 1.130 4.675 1.260 ;
        RECT 1.535 1.090 4.675 1.130 ;
        RECT 1.535 0.880 2.725 1.090 ;
        RECT 2.395 0.595 2.725 0.880 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.505 1.950 0.835 3.245 ;
        RECT 1.005 1.680 1.335 2.700 ;
        RECT 1.540 1.850 1.870 3.245 ;
        RECT 2.850 2.290 4.190 3.245 ;
        RECT 4.760 2.290 5.885 3.245 ;
        RECT 6.835 2.290 8.035 3.245 ;
        RECT 8.675 1.950 8.955 3.245 ;
        RECT 1.005 1.430 2.850 1.680 ;
        RECT 1.005 1.130 1.335 1.430 ;
        RECT 5.965 1.130 7.170 1.180 ;
        RECT 0.115 0.960 1.335 1.130 ;
        RECT 5.105 1.010 9.005 1.130 ;
        RECT 5.105 0.960 6.215 1.010 ;
        RECT 0.115 0.770 0.445 0.960 ;
        RECT 2.905 0.750 4.875 0.920 ;
        RECT 5.105 0.770 5.435 0.960 ;
        RECT 5.965 0.770 6.215 0.960 ;
        RECT 6.920 0.960 9.005 1.010 ;
        RECT 0.545 0.085 0.875 0.600 ;
        RECT 1.105 0.425 1.435 0.710 ;
        RECT 1.965 0.425 2.215 0.710 ;
        RECT 2.905 0.425 3.075 0.750 ;
        RECT 5.605 0.600 5.795 0.710 ;
        RECT 6.395 0.600 6.725 0.840 ;
        RECT 5.535 0.580 6.725 0.600 ;
        RECT 1.105 0.255 3.075 0.425 ;
        RECT 3.255 0.330 6.725 0.580 ;
        RECT 6.920 0.350 7.100 0.960 ;
        RECT 7.270 0.085 7.600 0.780 ;
        RECT 7.770 0.350 7.960 0.960 ;
        RECT 8.130 0.085 8.505 0.780 ;
        RECT 8.675 0.350 9.005 0.960 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__nand4b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.255 0.480 0.670 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.470 1.315 1.800 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.985 0.810 3.315 1.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 3.885 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 1.330 0.975 1.375 ;
        RECT 0.030 1.240 1.555 1.330 ;
        RECT 0.030 0.950 4.085 1.240 ;
        RECT 0.030 0.245 4.265 0.950 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.248650 ;
    PORT
      LAYER li1 ;
        RECT 1.675 2.480 2.005 2.980 ;
        RECT 2.765 2.480 3.095 2.980 ;
        RECT 1.675 2.310 3.095 2.480 ;
        RECT 2.525 2.120 3.095 2.310 ;
        RECT 3.765 2.120 4.225 2.980 ;
        RECT 2.525 1.950 4.225 2.120 ;
        RECT 2.525 1.820 3.095 1.950 ;
        RECT 4.055 1.180 4.225 1.950 ;
        RECT 3.485 1.010 4.225 1.180 ;
        RECT 3.485 0.620 3.655 1.010 ;
        RECT 1.720 0.350 3.655 0.620 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 1.970 0.445 2.850 ;
        RECT 0.615 1.970 0.945 3.245 ;
        RECT 1.115 2.140 1.445 2.850 ;
        RECT 2.175 2.650 2.595 3.245 ;
        RECT 3.265 2.290 3.595 3.245 ;
        RECT 1.115 1.970 2.355 2.140 ;
        RECT 0.115 1.300 0.285 1.970 ;
        RECT 2.185 1.550 2.355 1.970 ;
        RECT 1.685 1.300 2.015 1.550 ;
        RECT 0.115 1.130 2.015 1.300 ;
        RECT 2.185 1.220 2.745 1.550 ;
        RECT 0.115 0.840 0.470 1.130 ;
        RECT 2.185 0.960 2.355 1.220 ;
        RECT 0.650 0.085 0.980 0.960 ;
        RECT 1.150 0.790 2.355 0.960 ;
        RECT 1.150 0.630 1.490 0.790 ;
        RECT 3.825 0.085 4.155 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__nand4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.300 0.835 1.780 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.180 1.335 1.510 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 5.385 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.680 6.595 1.780 ;
        RECT 5.625 1.350 6.595 1.680 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.735 1.140 6.710 1.240 ;
        RECT 0.020 0.245 6.710 1.140 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.614500 ;
    PORT
      LAYER li1 ;
        RECT 2.345 2.020 2.675 2.980 ;
        RECT 3.345 2.120 3.675 2.980 ;
        RECT 4.775 2.120 5.105 2.980 ;
        RECT 5.775 2.120 6.105 2.980 ;
        RECT 3.345 2.020 6.105 2.120 ;
        RECT 2.345 1.950 6.105 2.020 ;
        RECT 2.345 1.850 4.195 1.950 ;
        RECT 5.775 1.850 6.105 1.950 ;
        RECT 2.345 1.820 2.675 1.850 ;
        RECT 3.965 1.260 4.195 1.850 ;
        RECT 2.685 1.090 4.195 1.260 ;
        RECT 2.685 0.840 2.855 1.090 ;
        RECT 2.345 0.670 2.855 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.095 2.410 0.445 2.860 ;
        RECT 0.650 2.580 0.980 3.245 ;
        RECT 1.845 2.580 2.175 3.245 ;
        RECT 0.095 2.240 2.175 2.410 ;
        RECT 0.095 1.950 0.445 2.240 ;
        RECT 0.095 1.030 0.265 1.950 ;
        RECT 1.185 1.820 1.675 2.070 ;
        RECT 1.505 1.180 1.675 1.820 ;
        RECT 1.845 1.350 2.175 2.240 ;
        RECT 2.845 2.190 3.175 3.245 ;
        RECT 3.845 2.290 4.605 3.245 ;
        RECT 5.275 2.290 5.605 3.245 ;
        RECT 6.275 1.950 6.605 3.245 ;
        RECT 3.125 1.600 3.795 1.680 ;
        RECT 2.345 1.430 3.795 1.600 ;
        RECT 2.345 1.180 2.515 1.430 ;
        RECT 0.095 0.350 0.460 1.030 ;
        RECT 1.505 1.010 2.515 1.180 ;
        RECT 4.410 1.010 6.600 1.180 ;
        RECT 0.630 0.085 0.960 1.010 ;
        RECT 1.130 0.350 1.675 1.010 ;
        RECT 1.845 0.500 2.175 0.840 ;
        RECT 3.025 0.750 4.180 0.920 ;
        RECT 3.025 0.500 3.195 0.750 ;
        RECT 4.410 0.620 4.740 1.010 ;
        RECT 1.845 0.330 3.195 0.500 ;
        RECT 3.365 0.425 3.695 0.580 ;
        RECT 4.910 0.425 5.240 0.815 ;
        RECT 3.365 0.255 5.240 0.425 ;
        RECT 5.420 0.350 5.670 1.010 ;
        RECT 5.840 0.085 6.170 0.815 ;
        RECT 6.350 0.350 6.600 1.010 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__nand4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 0.440 1.450 0.835 1.780 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.550 1.795 1.880 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.650 7.075 1.780 ;
        RECT 6.185 1.320 7.610 1.650 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.265 1.300 9.955 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 1.610 1.440 ;
        RECT 0.005 0.245 10.075 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.236100 ;
    PORT
      LAYER li1 ;
        RECT 2.525 2.230 2.965 2.990 ;
        RECT 3.635 2.230 3.865 2.990 ;
        RECT 4.535 2.230 4.815 2.980 ;
        RECT 2.525 2.060 4.815 2.230 ;
        RECT 4.485 2.020 4.815 2.060 ;
        RECT 5.515 2.020 5.685 2.980 ;
        RECT 4.485 1.990 5.685 2.020 ;
        RECT 6.335 2.120 6.665 2.980 ;
        RECT 7.335 2.120 7.665 2.980 ;
        RECT 8.285 2.120 8.615 2.980 ;
        RECT 9.185 2.120 9.515 2.980 ;
        RECT 6.335 1.990 9.515 2.120 ;
        RECT 4.485 1.950 9.515 1.990 ;
        RECT 4.485 1.850 6.665 1.950 ;
        RECT 5.515 1.820 6.665 1.850 ;
        RECT 7.335 1.820 7.665 1.950 ;
        RECT 5.515 1.260 5.685 1.820 ;
        RECT 3.335 1.090 5.685 1.260 ;
        RECT 3.335 1.040 3.505 1.090 ;
        RECT 2.320 0.870 3.505 1.040 ;
        RECT 2.320 0.595 2.650 0.870 ;
        RECT 3.335 0.595 3.505 0.870 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.115 2.290 0.445 3.245 ;
        RECT 0.645 2.120 0.815 2.980 ;
        RECT 1.015 2.390 1.345 3.245 ;
        RECT 1.515 2.220 1.795 2.980 ;
        RECT 2.005 2.390 2.335 3.245 ;
        RECT 3.135 2.400 3.465 3.245 ;
        RECT 4.035 2.400 4.365 3.245 ;
        RECT 0.100 1.950 0.815 2.120 ;
        RECT 1.125 2.050 2.135 2.220 ;
        RECT 4.985 2.190 5.315 3.245 ;
        RECT 5.885 2.160 6.135 3.245 ;
        RECT 6.835 2.290 7.165 3.245 ;
        RECT 7.865 2.290 8.115 3.245 ;
        RECT 8.815 2.290 8.985 3.245 ;
        RECT 0.100 1.280 0.270 1.950 ;
        RECT 1.125 1.330 1.295 2.050 ;
        RECT 1.965 1.890 2.135 2.050 ;
        RECT 9.715 1.950 9.965 3.245 ;
        RECT 1.965 1.720 4.315 1.890 ;
        RECT 4.145 1.680 4.315 1.720 ;
        RECT 2.155 1.380 3.165 1.550 ;
        RECT 4.145 1.430 5.345 1.680 ;
        RECT 0.100 0.830 0.445 1.280 ;
        RECT 1.125 1.000 1.420 1.330 ;
        RECT 1.590 1.210 3.165 1.380 ;
        RECT 1.590 0.830 1.760 1.210 ;
        RECT 6.125 1.130 8.095 1.150 ;
        RECT 0.100 0.660 1.760 0.830 ;
        RECT 0.100 0.550 0.445 0.660 ;
        RECT 0.625 0.085 0.955 0.490 ;
        RECT 1.930 0.425 2.100 1.040 ;
        RECT 6.125 0.980 9.965 1.130 ;
        RECT 3.685 0.750 5.895 0.920 ;
        RECT 2.820 0.425 3.150 0.700 ;
        RECT 3.685 0.425 3.935 0.750 ;
        RECT 5.565 0.595 5.895 0.750 ;
        RECT 6.125 0.595 6.375 0.980 ;
        RECT 1.930 0.255 3.935 0.425 ;
        RECT 4.115 0.425 5.385 0.580 ;
        RECT 6.555 0.425 6.885 0.810 ;
        RECT 7.065 0.595 7.235 0.980 ;
        RECT 7.925 0.960 9.965 0.980 ;
        RECT 7.415 0.425 7.745 0.810 ;
        RECT 4.115 0.255 7.745 0.425 ;
        RECT 7.925 0.350 8.095 0.960 ;
        RECT 8.275 0.085 8.605 0.790 ;
        RECT 8.785 0.350 8.955 0.960 ;
        RECT 9.135 0.085 9.465 0.790 ;
        RECT 9.635 0.350 9.965 0.960 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__nand4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.300 1.315 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 1.435 1.240 ;
        RECT 0.000 0.000 1.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.440 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.537600 ;
    PORT
      LAYER li1 ;
        RECT 0.985 2.890 1.315 2.980 ;
        RECT 0.645 1.950 1.315 2.890 ;
        RECT 0.645 1.130 0.815 1.950 ;
        RECT 0.565 0.350 0.815 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.440 3.415 ;
        RECT 0.115 1.950 0.445 3.245 ;
        RECT 0.135 0.085 0.385 1.130 ;
        RECT 0.995 0.085 1.325 1.130 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
  END
END sky130_fd_sc_hs__nor2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 1.410 2.135 1.605 ;
        RECT 1.805 0.440 2.275 1.410 ;
        RECT 1.805 0.255 2.135 0.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.180 0.445 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 1.555 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.820 0.945 2.735 ;
        RECT 0.615 0.350 0.945 1.820 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.155 2.905 1.305 3.075 ;
        RECT 0.155 1.820 0.405 2.905 ;
        RECT 1.135 1.945 1.305 2.905 ;
        RECT 1.505 2.115 1.755 3.245 ;
        RECT 1.955 1.945 2.285 2.980 ;
        RECT 1.135 1.775 2.285 1.945 ;
        RECT 0.115 0.085 0.445 1.010 ;
        RECT 1.115 0.085 1.445 1.130 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__nor2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 1.795 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.180 4.195 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.793600 ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.890 2.695 2.735 ;
        RECT 3.365 1.890 3.695 2.735 ;
        RECT 2.365 1.720 3.695 1.890 ;
        RECT 2.365 1.410 2.695 1.720 ;
        RECT 2.365 1.180 2.755 1.410 ;
        RECT 2.365 1.130 2.690 1.180 ;
        RECT 2.360 1.010 2.690 1.130 ;
        RECT 0.640 0.840 2.690 1.010 ;
        RECT 0.640 0.340 1.690 0.840 ;
        RECT 2.360 0.350 2.690 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 1.890 0.445 2.980 ;
        RECT 0.645 2.060 0.815 3.245 ;
        RECT 1.015 1.890 1.345 2.980 ;
        RECT 1.545 2.060 1.715 3.245 ;
        RECT 1.915 2.905 4.145 3.075 ;
        RECT 1.915 1.890 2.195 2.905 ;
        RECT 2.865 2.060 3.195 2.905 ;
        RECT 0.115 1.720 2.195 1.890 ;
        RECT 3.865 1.820 4.145 2.905 ;
        RECT 0.115 0.085 0.470 1.010 ;
        RECT 1.860 0.085 2.190 0.670 ;
        RECT 2.860 0.085 4.205 1.010 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__nor2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.788000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 3.715 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.788000 ;
    PORT
      LAYER li1 ;
        RECT 7.225 0.300 7.555 1.310 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.245 6.885 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.839300 ;
    PORT
      LAYER li1 ;
        RECT 4.415 1.780 4.745 2.735 ;
        RECT 5.365 1.780 5.695 2.735 ;
        RECT 4.415 1.650 5.695 1.780 ;
        RECT 6.265 1.650 6.595 2.735 ;
        RECT 7.215 1.650 7.545 2.735 ;
        RECT 4.415 1.480 7.545 1.650 ;
        RECT 4.415 1.310 6.275 1.480 ;
        RECT 4.260 1.180 6.275 1.310 ;
        RECT 1.860 1.140 6.275 1.180 ;
        RECT 1.860 1.010 5.275 1.140 ;
        RECT 1.860 0.350 2.190 1.010 ;
        RECT 3.260 0.350 3.590 1.010 ;
        RECT 4.260 0.350 5.275 1.010 ;
        RECT 5.945 0.350 6.275 1.140 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 1.950 0.445 2.980 ;
        RECT 0.615 2.120 0.945 3.245 ;
        RECT 1.145 2.120 1.315 2.980 ;
        RECT 1.515 2.290 1.845 3.245 ;
        RECT 2.045 2.120 2.295 2.980 ;
        RECT 2.465 2.290 2.795 3.245 ;
        RECT 2.995 2.120 3.245 2.980 ;
        RECT 3.415 2.290 3.745 3.245 ;
        RECT 3.915 2.905 8.045 3.075 ;
        RECT 3.915 2.120 4.245 2.905 ;
        RECT 1.145 1.950 4.245 2.120 ;
        RECT 4.925 1.950 5.185 2.905 ;
        RECT 0.115 1.780 1.315 1.950 ;
        RECT 5.875 1.820 6.080 2.905 ;
        RECT 6.775 1.820 7.035 2.905 ;
        RECT 7.715 1.820 8.045 2.905 ;
        RECT 0.650 0.085 1.690 1.130 ;
        RECT 2.360 0.085 3.090 0.840 ;
        RECT 3.760 0.085 4.090 0.840 ;
        RECT 5.445 0.085 5.775 0.970 ;
        RECT 6.445 0.085 6.775 1.130 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__nor2_8

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.180 1.365 1.550 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.180 0.440 1.550 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.682700 ;
    PORT
      LAYER li1 ;
        RECT 1.875 1.820 2.315 2.980 ;
        RECT 2.145 1.150 2.315 1.820 ;
        RECT 1.535 0.980 2.315 1.150 ;
        RECT 1.535 0.350 1.785 0.980 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.315 1.890 0.645 2.700 ;
        RECT 0.925 2.060 1.255 3.245 ;
        RECT 0.315 1.720 1.705 1.890 ;
        RECT 0.610 1.010 0.780 1.720 ;
        RECT 1.535 1.650 1.705 1.720 ;
        RECT 1.535 1.320 1.975 1.650 ;
        RECT 0.255 0.680 0.780 1.010 ;
        RECT 0.950 0.085 1.280 1.010 ;
        RECT 1.955 0.085 2.230 0.810 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__nor2b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.755 1.780 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.530 1.470 0.860 1.800 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.340 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824400 ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.180 1.820 2.735 ;
        RECT 3.005 1.180 3.235 1.410 ;
        RECT 1.645 1.010 3.235 1.180 ;
        RECT 1.645 0.960 2.745 1.010 ;
        RECT 1.485 0.350 1.815 0.960 ;
        RECT 2.495 0.350 2.745 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.110 1.300 0.360 2.980 ;
        RECT 0.560 1.970 0.890 3.245 ;
        RECT 1.120 2.905 2.350 3.075 ;
        RECT 1.120 1.820 1.450 2.905 ;
        RECT 2.020 2.120 2.350 2.905 ;
        RECT 2.550 2.290 2.800 3.245 ;
        RECT 3.000 2.120 3.250 2.980 ;
        RECT 2.020 1.950 3.250 2.120 ;
        RECT 3.000 1.820 3.250 1.950 ;
        RECT 1.145 1.300 1.475 1.550 ;
        RECT 0.110 1.130 1.475 1.300 ;
        RECT 0.110 0.450 0.780 1.130 ;
        RECT 0.985 0.085 1.315 0.960 ;
        RECT 1.985 0.085 2.315 0.790 ;
        RECT 2.915 0.085 3.245 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__nor2b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.340 1.795 1.410 ;
        RECT 0.790 1.180 1.795 1.340 ;
        RECT 3.645 1.180 3.975 1.550 ;
        RECT 0.790 1.010 3.975 1.180 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 4.750 1.180 5.155 1.825 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.440 0.245 5.275 1.240 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 1.885 2.230 2.165 2.735 ;
        RECT 2.895 2.230 3.145 2.735 ;
        RECT 1.885 2.060 3.145 2.230 ;
        RECT 1.885 1.850 2.165 2.060 ;
        RECT 1.885 1.750 2.055 1.850 ;
        RECT 0.535 1.680 2.055 1.750 ;
        RECT 0.185 1.580 2.055 1.680 ;
        RECT 0.185 1.510 0.705 1.580 ;
        RECT 0.185 1.410 0.355 1.510 ;
        RECT 0.125 0.840 0.355 1.410 ;
        RECT 0.125 0.670 3.810 0.840 ;
        RECT 2.060 0.530 2.390 0.670 ;
        RECT 3.560 0.510 3.810 0.670 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.115 1.850 0.365 3.245 ;
        RECT 0.565 2.090 0.895 2.980 ;
        RECT 1.095 2.260 1.265 3.245 ;
        RECT 1.465 2.905 3.645 3.075 ;
        RECT 1.465 2.090 1.715 2.905 ;
        RECT 2.365 2.400 2.695 2.905 ;
        RECT 0.565 1.920 1.715 2.090 ;
        RECT 3.315 2.060 3.645 2.905 ;
        RECT 3.815 2.060 4.145 3.245 ;
        RECT 4.350 1.995 4.680 2.875 ;
        RECT 4.880 1.995 5.130 3.245 ;
        RECT 4.350 1.890 4.580 1.995 ;
        RECT 3.055 1.720 4.580 1.890 ;
        RECT 3.055 1.680 3.225 1.720 ;
        RECT 2.225 1.350 3.225 1.680 ;
        RECT 4.410 1.010 4.580 1.720 ;
        RECT 1.550 0.085 1.880 0.500 ;
        RECT 2.570 0.085 3.380 0.500 ;
        RECT 3.990 0.085 4.240 0.840 ;
        RECT 4.410 0.345 5.165 1.010 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__nor2b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.360 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.870 1.300 1.315 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.300 1.815 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 1.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 1.915 1.240 ;
        RECT 0.000 0.000 1.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.110 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 1.920 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.737300 ;
    PORT
      LAYER li1 ;
        RECT 0.605 2.120 1.815 2.980 ;
        RECT 0.530 1.950 1.815 2.120 ;
        RECT 0.530 1.130 0.700 1.950 ;
        RECT 0.530 0.880 1.805 1.130 ;
        RECT 0.615 0.365 0.805 0.880 ;
        RECT 1.475 0.350 1.805 0.880 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 1.920 3.415 ;
        RECT 0.105 2.325 0.435 3.245 ;
        RECT 0.105 1.950 0.355 2.325 ;
        RECT 0.115 0.710 0.360 1.010 ;
        RECT 0.115 0.085 0.445 0.710 ;
        RECT 0.975 0.085 1.305 0.710 ;
        RECT 0.000 -0.085 1.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
  END
END sky130_fd_sc_hs__nor3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 2.650 0.310 3.235 0.980 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 1.305 1.380 3.255 1.550 ;
        RECT 1.305 1.220 1.635 1.380 ;
        RECT 2.925 1.180 3.255 1.380 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.180 0.975 1.550 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.590 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.861900 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.890 0.945 2.735 ;
        RECT 0.115 1.720 0.945 1.890 ;
        RECT 0.115 1.010 0.355 1.720 ;
        RECT 1.650 1.010 1.980 1.050 ;
        RECT 0.115 0.840 1.980 1.010 ;
        RECT 0.115 0.350 0.445 0.840 ;
        RECT 1.650 0.350 1.980 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.905 1.315 3.075 ;
        RECT 0.115 2.060 0.445 2.905 ;
        RECT 1.145 1.890 1.315 2.905 ;
        RECT 1.515 2.230 1.845 2.990 ;
        RECT 2.015 2.400 2.345 3.245 ;
        RECT 2.515 2.230 2.795 2.990 ;
        RECT 1.515 2.060 2.795 2.230 ;
        RECT 2.965 1.890 3.245 2.980 ;
        RECT 1.145 1.720 3.245 1.890 ;
        RECT 0.615 0.085 1.480 0.650 ;
        RECT 2.150 0.085 2.480 1.130 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__nor3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 1.625 2.190 4.020 2.340 ;
        RECT 1.625 2.170 6.135 2.190 ;
        RECT 0.605 1.920 1.795 2.170 ;
        RECT 3.850 2.020 6.135 2.170 ;
        RECT 0.605 1.350 0.935 1.920 ;
        RECT 5.805 0.330 6.135 2.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 1.310 1.520 1.640 1.680 ;
        RECT 1.310 1.510 2.755 1.520 ;
        RECT 1.310 1.350 4.965 1.510 ;
        RECT 2.045 1.180 4.965 1.350 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 3.785 0.340 5.635 0.670 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.670 1.240 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
        RECT 1.780 1.590 3.830 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.674800 ;
    PORT
      LAYER li1 ;
        RECT 2.140 1.850 3.680 2.000 ;
        RECT 2.140 1.750 5.305 1.850 ;
        RECT 3.350 1.680 5.305 1.750 ;
        RECT 0.545 1.010 1.875 1.180 ;
        RECT 5.135 1.010 5.305 1.680 ;
        RECT 0.545 0.350 0.875 1.010 ;
        RECT 1.545 0.840 5.305 1.010 ;
        RECT 1.545 0.350 1.875 0.840 ;
        RECT 2.545 0.350 2.875 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.110 2.510 0.360 2.980 ;
        RECT 0.560 2.680 0.890 3.245 ;
        RECT 1.090 2.680 1.340 2.980 ;
        RECT 1.540 2.905 5.265 3.075 ;
        RECT 1.540 2.850 4.285 2.905 ;
        RECT 4.485 2.680 4.735 2.735 ;
        RECT 4.935 2.700 5.265 2.905 ;
        RECT 1.090 2.530 4.735 2.680 ;
        RECT 5.465 2.530 5.635 3.000 ;
        RECT 5.835 2.700 6.165 3.245 ;
        RECT 6.365 2.530 6.615 2.980 ;
        RECT 1.090 2.510 6.615 2.530 ;
        RECT 0.110 2.340 1.340 2.510 ;
        RECT 4.485 2.360 6.615 2.510 ;
        RECT 0.110 1.820 0.360 2.340 ;
        RECT 6.365 1.820 6.615 2.360 ;
        RECT 0.115 0.085 0.365 1.130 ;
        RECT 1.045 0.085 1.375 0.840 ;
        RECT 2.045 0.085 2.375 0.670 ;
        RECT 3.055 0.085 3.365 0.670 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__nor3_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.350 1.315 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.555 1.350 1.885 1.780 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.180 0.815 1.550 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.770 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.778100 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.290 2.795 2.980 ;
        RECT 2.625 1.180 2.795 2.290 ;
        RECT 1.330 1.010 2.795 1.180 ;
        RECT 1.330 0.350 1.660 1.010 ;
        RECT 2.330 0.350 2.795 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.105 2.120 0.595 2.700 ;
        RECT 0.835 2.290 1.165 3.245 ;
        RECT 0.105 1.950 2.295 2.120 ;
        RECT 0.105 1.820 0.595 1.950 ;
        RECT 0.105 1.010 0.275 1.820 ;
        RECT 2.125 1.680 2.295 1.950 ;
        RECT 2.125 1.350 2.455 1.680 ;
        RECT 0.105 0.680 0.650 1.010 ;
        RECT 0.830 0.085 1.160 1.010 ;
        RECT 1.830 0.085 2.160 0.840 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__nor3b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.675 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.605 1.350 3.275 1.780 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.450 0.835 1.780 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.615 1.140 4.795 1.240 ;
        RECT 0.010 0.245 4.795 1.140 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.005700 ;
    PORT
      LAYER li1 ;
        RECT 1.640 1.130 1.810 2.735 ;
        RECT 1.565 0.960 4.185 1.130 ;
        RECT 1.565 0.940 2.695 0.960 ;
        RECT 1.120 0.770 2.695 0.940 ;
        RECT 1.120 0.350 1.395 0.770 ;
        RECT 2.505 0.350 2.695 0.770 ;
        RECT 3.925 0.350 4.185 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.085 1.950 0.360 2.980 ;
        RECT 0.560 1.950 0.890 3.245 ;
        RECT 1.110 2.905 3.240 3.075 ;
        RECT 0.085 1.280 0.255 1.950 ;
        RECT 1.110 1.820 1.440 2.905 ;
        RECT 2.010 1.820 2.290 2.905 ;
        RECT 2.460 2.120 2.790 2.735 ;
        RECT 2.970 2.290 3.240 2.905 ;
        RECT 3.460 2.290 3.790 3.245 ;
        RECT 3.990 2.120 4.240 2.980 ;
        RECT 2.460 1.950 4.240 2.120 ;
        RECT 4.425 1.950 4.690 3.245 ;
        RECT 1.005 1.280 1.335 1.550 ;
        RECT 0.085 1.110 1.335 1.280 ;
        RECT 0.085 0.350 0.450 1.110 ;
        RECT 0.620 0.085 0.950 0.940 ;
        RECT 1.565 0.085 2.335 0.600 ;
        RECT 2.865 0.085 3.755 0.770 ;
        RECT 4.355 0.085 4.685 1.130 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__nor3b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.440 1.220 6.595 1.550 ;
        RECT 6.365 1.180 6.595 1.220 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.815 1.780 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.180 7.095 1.550 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 7.675 1.240 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.985500 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.820 3.720 2.070 ;
        RECT 2.045 1.180 2.275 1.820 ;
        RECT 0.615 1.150 2.275 1.180 ;
        RECT 0.615 1.050 3.805 1.150 ;
        RECT 0.615 1.010 5.935 1.050 ;
        RECT 0.615 0.350 0.945 1.010 ;
        RECT 1.615 0.980 5.935 1.010 ;
        RECT 1.615 0.350 1.945 0.980 ;
        RECT 2.625 0.350 2.795 0.980 ;
        RECT 3.475 0.880 5.935 0.980 ;
        RECT 3.475 0.350 3.805 0.880 ;
        RECT 4.475 0.350 4.805 0.880 ;
        RECT 5.605 0.350 5.935 0.880 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.115 2.905 2.370 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 0.615 2.120 0.945 2.735 ;
        RECT 1.145 2.290 1.315 2.905 ;
        RECT 2.040 2.750 2.370 2.905 ;
        RECT 2.940 2.750 3.270 2.910 ;
        RECT 3.840 2.750 4.170 2.910 ;
        RECT 1.525 2.410 1.855 2.735 ;
        RECT 2.040 2.580 4.170 2.750 ;
        RECT 4.400 2.580 4.730 3.245 ;
        RECT 4.930 2.410 5.100 2.990 ;
        RECT 1.525 2.240 5.100 2.410 ;
        RECT 5.300 2.400 5.630 3.245 ;
        RECT 1.525 2.120 1.870 2.240 ;
        RECT 0.615 1.950 1.870 2.120 ;
        RECT 4.795 2.230 5.100 2.240 ;
        RECT 5.810 2.230 6.080 2.990 ;
        RECT 4.795 2.060 6.080 2.230 ;
        RECT 6.250 2.060 6.580 3.245 ;
        RECT 6.785 1.890 7.055 2.700 ;
        RECT 7.235 2.060 7.565 3.245 ;
        RECT 3.890 1.720 7.565 1.890 ;
        RECT 3.890 1.650 4.195 1.720 ;
        RECT 2.580 1.320 4.195 1.650 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 7.395 1.010 7.565 1.720 ;
        RECT 1.115 0.085 1.445 0.840 ;
        RECT 2.115 0.085 2.445 0.810 ;
        RECT 2.975 0.085 3.305 0.810 ;
        RECT 3.975 0.085 4.305 0.710 ;
        RECT 4.975 0.085 5.435 0.680 ;
        RECT 6.105 0.085 6.435 1.010 ;
        RECT 6.605 0.350 7.565 1.010 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__nor3b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.540 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.350 1.315 2.890 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 2.150 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.445 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.950 2.645 1.240 ;
        RECT 0.100 0.245 2.750 0.950 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.744800 ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.950 2.785 2.980 ;
        RECT 2.615 1.180 2.785 1.950 ;
        RECT 0.780 1.010 2.785 1.180 ;
        RECT 0.780 0.350 1.040 1.010 ;
        RECT 1.810 0.350 2.140 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.255 1.820 0.585 3.245 ;
        RECT 0.210 0.085 0.610 1.010 ;
        RECT 1.210 0.085 1.540 0.840 ;
        RECT 2.310 0.085 2.640 0.840 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__nor4_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.180 3.715 1.540 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 2.455 1.710 4.215 1.880 ;
        RECT 2.455 1.650 2.625 1.710 ;
        RECT 2.285 1.320 2.625 1.650 ;
        RECT 3.885 0.280 4.215 1.710 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.650 1.795 2.150 ;
        RECT 1.565 1.500 2.075 1.650 ;
        RECT 0.425 1.320 2.075 1.500 ;
        RECT 0.425 1.170 0.700 1.320 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.330 0.435 0.660 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.005 0.790 3.490 1.240 ;
        RECT 0.495 0.245 3.490 0.790 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.808000 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.840 1.385 2.150 ;
        RECT 0.085 1.670 1.385 1.840 ;
        RECT 0.085 1.000 0.255 1.670 ;
        RECT 1.550 1.000 2.880 1.150 ;
        RECT 0.085 0.980 2.880 1.000 ;
        RECT 0.085 0.830 1.880 0.980 ;
        RECT 1.550 0.350 1.880 0.830 ;
        RECT 2.550 0.350 2.880 0.980 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.490 0.365 3.000 ;
        RECT 0.565 2.660 1.835 2.980 ;
        RECT 2.035 2.490 2.285 2.980 ;
        RECT 0.115 2.320 2.285 2.490 ;
        RECT 2.475 2.560 2.805 3.000 ;
        RECT 2.975 2.730 3.305 3.245 ;
        RECT 3.505 2.560 3.755 3.000 ;
        RECT 2.475 2.390 3.755 2.560 ;
        RECT 0.115 2.010 0.445 2.320 ;
        RECT 2.035 2.220 2.285 2.320 ;
        RECT 3.940 2.220 4.205 2.980 ;
        RECT 2.035 2.050 4.205 2.220 ;
        RECT 2.035 1.820 2.285 2.050 ;
        RECT 0.605 0.085 1.380 0.600 ;
        RECT 2.050 0.085 2.380 0.810 ;
        RECT 3.050 0.085 3.380 1.010 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__nor4_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 7.045 1.300 8.515 1.630 ;
        RECT 7.805 1.180 8.515 1.300 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 6.595 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.350 3.785 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.894000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.350 1.875 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 8.470 1.240 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.214400 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.120 0.945 2.735 ;
        RECT 1.565 2.120 1.895 2.735 ;
        RECT 0.125 1.950 1.895 2.120 ;
        RECT 0.125 1.180 0.355 1.950 ;
        RECT 0.125 1.130 4.590 1.180 ;
        RECT 0.125 1.010 7.570 1.130 ;
        RECT 0.615 0.350 1.740 1.010 ;
        RECT 2.410 0.350 3.590 1.010 ;
        RECT 4.260 0.960 7.860 1.010 ;
        RECT 4.260 0.350 4.590 0.960 ;
        RECT 7.240 0.340 7.860 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.115 2.905 2.265 3.075 ;
        RECT 0.115 2.290 0.445 2.905 ;
        RECT 1.145 2.290 1.395 2.905 ;
        RECT 2.095 2.120 2.265 2.905 ;
        RECT 2.465 2.905 6.075 3.075 ;
        RECT 2.465 2.290 2.795 2.905 ;
        RECT 2.970 2.120 3.190 2.735 ;
        RECT 3.365 2.290 3.695 2.905 ;
        RECT 3.895 2.120 4.145 2.735 ;
        RECT 2.095 1.950 4.145 2.120 ;
        RECT 4.375 2.120 4.625 2.735 ;
        RECT 4.825 2.300 5.155 2.905 ;
        RECT 5.340 2.120 5.560 2.735 ;
        RECT 5.745 2.300 6.075 2.905 ;
        RECT 6.255 2.120 6.525 2.980 ;
        RECT 6.695 2.290 7.025 3.245 ;
        RECT 7.195 2.120 7.525 2.980 ;
        RECT 7.695 2.290 8.025 3.245 ;
        RECT 8.195 2.120 8.525 2.980 ;
        RECT 4.375 1.950 8.525 2.120 ;
        RECT 2.095 1.820 2.265 1.950 ;
        RECT 8.195 1.820 8.525 1.950 ;
        RECT 0.115 0.085 0.445 0.840 ;
        RECT 1.910 0.085 2.240 0.840 ;
        RECT 3.760 0.085 4.090 0.840 ;
        RECT 4.760 0.085 7.070 0.790 ;
        RECT 8.030 0.085 8.360 1.010 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__nor4_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.350 1.315 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.350 1.855 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.395 1.780 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.110 0.815 1.440 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.785 1.050 3.240 1.240 ;
        RECT 0.180 0.245 3.240 1.050 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.879200 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.850 3.275 2.980 ;
        RECT 3.105 1.180 3.275 1.850 ;
        RECT 1.290 1.010 3.275 1.180 ;
        RECT 1.290 0.350 1.620 1.010 ;
        RECT 2.300 0.350 2.630 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.105 2.120 0.595 2.700 ;
        RECT 0.835 2.290 1.165 3.245 ;
        RECT 0.105 1.950 2.735 2.120 ;
        RECT 0.105 1.820 0.595 1.950 ;
        RECT 0.105 0.940 0.275 1.820 ;
        RECT 2.565 1.680 2.735 1.950 ;
        RECT 2.565 1.350 2.935 1.680 ;
        RECT 0.105 0.350 0.620 0.940 ;
        RECT 0.790 0.085 1.120 0.940 ;
        RECT 1.790 0.085 2.120 0.840 ;
        RECT 2.800 0.085 3.130 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__nor4b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 5.635 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.295 1.350 4.195 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.755 1.780 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.470 0.865 1.800 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.745 1.140 5.755 1.240 ;
        RECT 0.140 0.245 5.755 1.140 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.323900 ;
    PORT
      LAYER li1 ;
        RECT 1.655 2.120 1.825 2.735 ;
        RECT 1.655 1.950 3.095 2.120 ;
        RECT 1.655 1.820 1.825 1.950 ;
        RECT 2.925 1.180 3.095 1.950 ;
        RECT 2.440 1.010 5.145 1.180 ;
        RECT 2.440 0.960 2.770 1.010 ;
        RECT 1.250 0.790 2.770 0.960 ;
        RECT 1.250 0.330 1.580 0.790 ;
        RECT 2.440 0.350 2.770 0.790 ;
        RECT 3.440 0.350 3.770 1.010 ;
        RECT 4.815 0.350 5.145 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 1.300 0.365 2.980 ;
        RECT 0.565 1.970 0.895 3.245 ;
        RECT 1.125 2.905 2.275 3.075 ;
        RECT 1.125 1.820 1.455 2.905 ;
        RECT 2.025 2.460 2.275 2.905 ;
        RECT 2.475 2.905 4.265 3.075 ;
        RECT 2.475 2.630 2.805 2.905 ;
        RECT 3.005 2.460 3.255 2.735 ;
        RECT 2.025 2.290 3.255 2.460 ;
        RECT 3.485 2.120 3.735 2.735 ;
        RECT 3.935 2.290 4.265 2.905 ;
        RECT 4.465 2.120 4.635 2.980 ;
        RECT 4.835 2.290 5.165 3.245 ;
        RECT 5.375 2.120 5.625 2.980 ;
        RECT 3.485 1.950 5.625 2.120 ;
        RECT 1.105 1.300 1.775 1.550 ;
        RECT 0.115 1.130 1.775 1.300 ;
        RECT 0.115 0.350 0.580 1.130 ;
        RECT 0.750 0.085 1.080 0.960 ;
        RECT 1.750 0.085 2.270 0.600 ;
        RECT 2.940 0.085 3.270 0.840 ;
        RECT 3.940 0.085 4.645 0.790 ;
        RECT 5.315 0.085 5.645 1.130 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__nor4b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.350 9.475 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.350 7.555 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 3.920 1.350 5.155 1.780 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.920 0.550 1.930 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.540 0.860 10.075 1.240 ;
        RECT 0.105 0.245 10.075 0.860 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.440600 ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.990 2.355 2.735 ;
        RECT 2.975 2.120 3.305 2.735 ;
        RECT 2.975 1.990 5.635 2.120 ;
        RECT 2.025 1.950 5.635 1.990 ;
        RECT 2.025 1.820 3.305 1.950 ;
        RECT 2.500 1.300 3.750 1.470 ;
        RECT 2.500 1.150 2.830 1.300 ;
        RECT 1.570 0.980 2.830 1.150 ;
        RECT 1.570 0.350 1.820 0.980 ;
        RECT 2.500 0.350 2.830 0.980 ;
        RECT 3.500 1.180 3.750 1.300 ;
        RECT 5.405 1.180 5.635 1.950 ;
        RECT 3.500 1.010 9.465 1.180 ;
        RECT 3.500 0.350 3.750 1.010 ;
        RECT 4.905 0.350 5.235 1.010 ;
        RECT 6.250 0.350 6.580 1.010 ;
        RECT 7.250 0.350 7.580 1.010 ;
        RECT 8.275 0.350 8.525 1.010 ;
        RECT 9.215 0.350 9.465 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.115 2.100 0.365 3.245 ;
        RECT 0.565 2.100 0.895 2.980 ;
        RECT 1.075 2.100 1.345 3.245 ;
        RECT 1.575 2.905 3.755 3.075 ;
        RECT 0.720 1.650 0.890 2.100 ;
        RECT 1.575 1.820 1.825 2.905 ;
        RECT 2.525 2.160 2.805 2.905 ;
        RECT 3.475 2.490 3.755 2.905 ;
        RECT 3.925 2.905 7.715 3.075 ;
        RECT 3.925 2.660 4.255 2.905 ;
        RECT 4.425 2.490 4.755 2.720 ;
        RECT 4.925 2.630 5.255 2.905 ;
        RECT 3.475 2.460 4.755 2.490 ;
        RECT 5.440 2.460 5.705 2.540 ;
        RECT 3.475 2.320 5.705 2.460 ;
        RECT 4.425 2.290 5.705 2.320 ;
        RECT 5.935 2.120 6.265 2.735 ;
        RECT 6.435 2.290 6.765 2.905 ;
        RECT 6.935 2.120 7.265 2.735 ;
        RECT 7.465 2.290 7.715 2.905 ;
        RECT 7.885 2.120 8.115 2.980 ;
        RECT 8.285 2.290 8.535 3.245 ;
        RECT 8.735 2.120 9.065 2.980 ;
        RECT 9.265 2.290 9.515 3.245 ;
        RECT 9.715 2.120 9.965 2.980 ;
        RECT 5.935 1.950 9.965 2.120 ;
        RECT 9.715 1.820 9.965 1.950 ;
        RECT 0.720 1.320 2.330 1.650 ;
        RECT 0.720 0.750 0.890 1.320 ;
        RECT 0.275 0.420 0.890 0.750 ;
        RECT 1.060 0.085 1.390 1.130 ;
        RECT 2.000 0.085 2.330 0.790 ;
        RECT 3.000 0.085 3.330 1.130 ;
        RECT 3.930 0.085 4.735 0.840 ;
        RECT 5.405 0.085 6.080 0.840 ;
        RECT 6.750 0.085 7.080 0.805 ;
        RECT 7.750 0.085 8.105 0.805 ;
        RECT 8.705 0.085 9.035 0.805 ;
        RECT 9.635 0.085 9.965 1.130 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__nor4b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.075 1.350 1.405 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.915 1.350 2.275 1.780 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.450 4.345 1.780 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.848400 ;
    PORT
      LAYER li1 ;
        RECT 1.575 2.060 3.455 2.390 ;
        RECT 1.575 1.130 1.745 2.060 ;
        RECT 1.445 1.050 1.775 1.130 ;
        RECT 1.445 0.880 3.235 1.050 ;
        RECT 1.445 0.350 1.775 0.880 ;
        RECT 2.860 0.350 3.235 0.880 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.650 2.900 1.345 3.245 ;
        RECT 0.115 2.560 3.795 2.730 ;
        RECT 0.115 1.820 0.775 2.560 ;
        RECT 3.625 1.890 3.795 2.560 ;
        RECT 3.965 2.100 4.185 3.245 ;
        RECT 4.355 2.100 4.685 2.980 ;
        RECT 0.605 1.010 0.775 1.820 ;
        RECT 2.485 1.720 3.795 1.890 ;
        RECT 2.485 1.350 2.815 1.720 ;
        RECT 3.070 1.260 3.740 1.550 ;
        RECT 4.515 1.260 4.685 2.100 ;
        RECT 3.070 1.220 4.685 1.260 ;
        RECT 0.115 0.680 0.775 1.010 ;
        RECT 0.945 0.085 1.275 1.130 ;
        RECT 3.570 1.090 4.685 1.220 ;
        RECT 1.945 0.085 2.690 0.680 ;
        RECT 3.405 0.085 4.175 0.920 ;
        RECT 4.355 0.540 4.685 1.090 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__nor4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 6.310 1.350 7.075 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.635 6.115 1.780 ;
        RECT 4.860 1.350 6.115 1.635 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.470 1.315 1.800 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.470 1.825 1.800 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.240 2.075 1.390 ;
        RECT 0.995 1.140 7.195 1.240 ;
        RECT 0.375 0.245 7.195 1.140 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.198100 ;
    PORT
      LAYER li1 ;
        RECT 2.975 2.020 3.225 2.735 ;
        RECT 2.975 1.850 4.285 2.020 ;
        RECT 4.115 1.780 4.285 1.850 ;
        RECT 4.115 1.550 4.675 1.780 ;
        RECT 4.115 1.180 4.285 1.550 ;
        RECT 3.955 1.010 6.575 1.180 ;
        RECT 3.955 0.840 4.285 1.010 ;
        RECT 2.890 0.670 4.285 0.840 ;
        RECT 2.890 0.350 3.220 0.670 ;
        RECT 3.955 0.350 4.285 0.670 ;
        RECT 4.965 0.350 5.215 1.010 ;
        RECT 6.325 0.350 6.575 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.115 1.970 0.445 2.980 ;
        RECT 0.615 1.970 1.715 3.245 ;
        RECT 1.885 2.140 2.215 2.980 ;
        RECT 2.495 2.905 3.725 3.075 ;
        RECT 1.885 1.970 2.325 2.140 ;
        RECT 0.115 1.300 0.285 1.970 ;
        RECT 2.155 1.680 2.325 1.970 ;
        RECT 2.495 1.850 2.775 2.905 ;
        RECT 3.395 2.360 3.725 2.905 ;
        RECT 3.895 2.905 5.685 3.075 ;
        RECT 3.895 2.530 4.175 2.905 ;
        RECT 4.345 2.360 4.675 2.735 ;
        RECT 3.395 2.190 4.675 2.360 ;
        RECT 4.905 2.120 5.155 2.735 ;
        RECT 5.355 2.290 5.685 2.905 ;
        RECT 5.855 2.120 6.185 2.980 ;
        RECT 6.385 2.290 6.555 3.245 ;
        RECT 6.755 2.120 7.085 2.980 ;
        RECT 4.905 1.950 7.085 2.120 ;
        RECT 4.905 1.820 5.155 1.950 ;
        RECT 2.155 1.350 3.165 1.680 ;
        RECT 3.615 1.350 3.945 1.680 ;
        RECT 2.155 1.300 2.325 1.350 ;
        RECT 0.115 1.130 0.815 1.300 ;
        RECT 0.485 0.880 0.815 1.130 ;
        RECT 1.620 1.050 2.325 1.300 ;
        RECT 3.615 1.180 3.785 1.350 ;
        RECT 2.495 1.010 3.785 1.180 ;
        RECT 2.495 0.880 2.665 1.010 ;
        RECT 0.485 0.710 2.665 0.880 ;
        RECT 0.485 0.360 0.815 0.710 ;
        RECT 0.990 0.085 1.515 0.540 ;
        RECT 2.195 0.085 2.710 0.540 ;
        RECT 3.400 0.085 3.775 0.500 ;
        RECT 4.455 0.085 4.785 0.840 ;
        RECT 5.385 0.085 6.155 0.840 ;
        RECT 6.755 0.085 7.085 1.130 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__nor4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hs__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.180 2.495 1.540 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.710 2.890 1.880 ;
        RECT 1.085 1.650 1.315 1.710 ;
        RECT 0.265 1.320 1.315 1.650 ;
        RECT 2.720 1.585 2.890 1.710 ;
        RECT 2.720 1.255 3.920 1.585 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 9.095 1.530 9.955 1.860 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 10.125 1.450 10.455 1.780 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 11.035 1.240 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
        RECT 2.480 1.565 8.675 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.544200 ;
    PORT
      LAYER li1 ;
        RECT 5.990 1.725 7.230 2.055 ;
        RECT 5.990 1.470 6.320 1.725 ;
        RECT 5.525 1.300 6.615 1.470 ;
        RECT 0.615 1.010 0.945 1.130 ;
        RECT 5.525 1.085 5.775 1.300 ;
        RECT 2.665 1.010 5.775 1.085 ;
        RECT 0.615 0.915 5.775 1.010 ;
        RECT 0.615 0.840 2.915 0.915 ;
        RECT 0.615 0.350 0.945 0.840 ;
        RECT 1.615 0.350 1.945 0.840 ;
        RECT 2.665 0.350 2.915 0.840 ;
        RECT 3.595 0.350 3.845 0.915 ;
        RECT 4.515 0.350 4.845 0.915 ;
        RECT 5.525 0.350 5.775 0.915 ;
        RECT 6.445 1.055 6.615 1.300 ;
        RECT 6.445 0.885 8.035 1.055 ;
        RECT 6.445 0.350 6.775 0.885 ;
        RECT 7.705 0.350 8.035 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.115 2.220 0.445 2.980 ;
        RECT 0.615 2.560 0.945 2.980 ;
        RECT 1.115 2.730 1.445 3.245 ;
        RECT 1.645 2.560 1.895 2.980 ;
        RECT 2.065 2.730 2.435 3.245 ;
        RECT 2.635 2.905 3.890 3.075 ;
        RECT 2.635 2.560 2.885 2.905 ;
        RECT 0.615 2.390 2.885 2.560 ;
        RECT 3.060 2.220 3.390 2.735 ;
        RECT 0.115 2.050 3.390 2.220 ;
        RECT 3.560 2.095 3.890 2.905 ;
        RECT 4.090 2.905 8.490 3.075 ;
        RECT 0.115 1.820 0.445 2.050 ;
        RECT 3.060 1.925 3.390 2.050 ;
        RECT 4.090 1.925 4.260 2.905 ;
        RECT 3.060 1.755 4.260 1.925 ;
        RECT 4.470 2.565 8.035 2.735 ;
        RECT 4.470 1.755 4.800 2.565 ;
        RECT 5.185 2.225 7.570 2.395 ;
        RECT 5.185 1.585 5.355 2.225 ;
        RECT 7.400 1.895 7.570 2.225 ;
        RECT 7.760 2.065 8.035 2.565 ;
        RECT 8.205 2.065 8.490 2.905 ;
        RECT 8.790 2.370 9.120 3.245 ;
        RECT 9.300 2.200 9.575 2.980 ;
        RECT 8.705 2.030 9.575 2.200 ;
        RECT 9.775 2.100 9.945 3.245 ;
        RECT 10.145 2.120 10.395 2.980 ;
        RECT 10.595 2.290 10.925 3.245 ;
        RECT 8.705 1.895 8.875 2.030 ;
        RECT 10.145 1.950 10.925 2.120 ;
        RECT 7.400 1.725 8.875 1.895 ;
        RECT 4.345 1.255 5.355 1.585 ;
        RECT 6.785 1.225 8.375 1.555 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 1.115 0.085 1.445 0.670 ;
        RECT 2.115 0.085 2.445 0.670 ;
        RECT 3.085 0.085 3.415 0.745 ;
        RECT 4.015 0.085 4.345 0.745 ;
        RECT 5.015 0.085 5.345 0.745 ;
        RECT 5.945 0.085 6.275 1.130 ;
        RECT 8.205 1.020 8.375 1.225 ;
        RECT 8.545 1.360 8.875 1.725 ;
        RECT 8.545 1.190 9.585 1.360 ;
        RECT 10.755 1.280 10.925 1.950 ;
        RECT 8.205 0.850 9.090 1.020 ;
        RECT 6.945 0.085 7.535 0.680 ;
        RECT 8.205 0.085 8.750 0.680 ;
        RECT 8.920 0.425 9.090 0.850 ;
        RECT 9.260 0.670 9.585 1.190 ;
        RECT 9.755 1.110 10.925 1.280 ;
        RECT 9.755 0.425 9.925 1.110 ;
        RECT 8.920 0.255 9.925 0.425 ;
        RECT 10.095 0.085 10.495 0.940 ;
        RECT 10.665 0.350 10.925 1.110 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__nor4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2bb2a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.710 1.315 1.780 ;
        RECT 0.965 1.420 1.315 1.710 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.430 1.835 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.180 4.215 1.510 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.180 3.715 1.510 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 1.140 2.070 1.240 ;
        RECT 0.015 0.245 4.315 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.445 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.455 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.615 1.950 0.945 3.245 ;
        RECT 1.655 2.450 2.820 3.245 ;
        RECT 1.150 1.950 2.380 2.280 ;
        RECT 2.990 2.070 3.320 2.780 ;
        RECT 0.425 1.300 0.795 1.630 ;
        RECT 0.625 1.250 0.795 1.300 ;
        RECT 2.050 1.260 2.380 1.950 ;
        RECT 0.625 1.080 1.460 1.250 ;
        RECT 0.625 0.085 1.120 0.910 ;
        RECT 1.290 0.425 1.460 1.080 ;
        RECT 1.630 1.090 2.380 1.260 ;
        RECT 2.645 1.900 3.320 2.070 ;
        RECT 3.870 1.900 4.200 3.245 ;
        RECT 1.630 0.595 1.880 1.090 ;
        RECT 2.645 0.920 2.815 1.900 ;
        RECT 2.485 0.425 2.815 0.920 ;
        RECT 1.290 0.255 2.815 0.425 ;
        RECT 2.995 0.840 4.205 1.010 ;
        RECT 2.995 0.340 3.245 0.840 ;
        RECT 3.415 0.085 3.745 0.670 ;
        RECT 3.955 0.340 4.205 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o2bb2a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o2bb2a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2bb2a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.475 2.865 1.805 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.475 2.325 1.805 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.570 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.810 1.450 1.285 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 1.915 1.240 ;
        RECT 2.925 1.140 4.300 1.240 ;
        RECT 0.005 0.245 4.300 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.425 1.820 3.770 2.980 ;
        RECT 3.600 1.130 3.770 1.820 ;
        RECT 3.430 0.350 3.770 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.120 1.950 0.450 3.245 ;
        RECT 1.050 2.565 1.380 2.980 ;
        RECT 1.585 2.735 1.940 3.245 ;
        RECT 2.770 2.735 3.220 3.245 ;
        RECT 1.050 2.395 3.255 2.565 ;
        RECT 1.050 1.950 1.380 2.395 ;
        RECT 1.615 1.975 2.565 2.225 ;
        RECT 1.615 1.780 1.785 1.975 ;
        RECT 1.455 1.450 1.785 1.780 ;
        RECT 1.615 1.305 1.785 1.450 ;
        RECT 3.085 1.635 3.255 2.395 ;
        RECT 3.955 1.820 4.205 3.245 ;
        RECT 3.085 1.305 3.430 1.635 ;
        RECT 0.115 1.110 1.305 1.280 ;
        RECT 1.615 1.135 2.375 1.305 ;
        RECT 0.115 0.350 0.365 1.110 ;
        RECT 0.545 0.085 0.875 0.940 ;
        RECT 1.055 0.350 1.305 1.110 ;
        RECT 1.475 0.425 1.805 0.965 ;
        RECT 2.045 0.595 2.375 1.135 ;
        RECT 2.545 1.135 3.255 1.305 ;
        RECT 2.545 0.425 2.715 1.135 ;
        RECT 1.475 0.255 2.715 0.425 ;
        RECT 2.885 0.085 3.215 0.965 ;
        RECT 3.940 0.085 4.190 1.130 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o2bb2a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2bb2a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 4.415 1.350 4.745 1.780 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 3.845 1.350 4.195 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.260 1.115 1.770 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.470 1.450 2.275 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.590 1.140 7.195 1.240 ;
        RECT 0.005 0.245 7.195 1.140 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.311300 ;
    PORT
      LAYER li1 ;
        RECT 5.255 1.890 5.585 2.980 ;
        RECT 6.255 1.890 6.585 2.980 ;
        RECT 5.255 1.720 6.585 1.890 ;
        RECT 6.255 1.050 6.585 1.720 ;
        RECT 5.255 0.810 6.585 1.050 ;
        RECT 5.255 0.350 5.585 0.810 ;
        RECT 6.255 0.350 6.585 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.185 2.120 0.515 2.980 ;
        RECT 0.715 2.290 0.885 3.245 ;
        RECT 1.085 2.905 2.315 3.075 ;
        RECT 1.085 2.120 1.415 2.905 ;
        RECT 0.185 1.950 1.415 2.120 ;
        RECT 1.615 2.120 1.785 2.735 ;
        RECT 1.985 2.290 2.315 2.905 ;
        RECT 2.545 2.320 2.875 3.245 ;
        RECT 3.600 2.790 3.930 3.245 ;
        RECT 4.670 2.790 5.000 3.245 ;
        RECT 3.165 2.450 5.085 2.620 ;
        RECT 3.165 2.150 3.335 2.450 ;
        RECT 2.995 2.120 3.335 2.150 ;
        RECT 1.615 1.950 3.335 2.120 ;
        RECT 0.185 1.940 0.515 1.950 ;
        RECT 2.995 1.820 3.335 1.950 ;
        RECT 3.505 1.950 4.465 2.280 ;
        RECT 3.505 1.630 3.675 1.950 ;
        RECT 2.490 1.300 3.675 1.630 ;
        RECT 3.505 1.130 3.675 1.300 ;
        RECT 4.915 1.550 5.085 2.450 ;
        RECT 5.755 2.060 6.085 3.245 ;
        RECT 6.755 1.820 7.085 3.245 ;
        RECT 4.915 1.220 6.065 1.550 ;
        RECT 0.115 0.920 3.335 1.090 ;
        RECT 3.505 0.960 4.030 1.130 ;
        RECT 4.915 1.120 5.085 1.220 ;
        RECT 0.115 0.350 0.445 0.920 ;
        RECT 1.115 0.780 3.335 0.920 ;
        RECT 0.615 0.085 0.945 0.750 ;
        RECT 1.115 0.350 1.445 0.780 ;
        RECT 1.615 0.085 1.945 0.610 ;
        RECT 2.505 0.425 2.835 0.610 ;
        RECT 3.005 0.595 3.335 0.780 ;
        RECT 3.700 0.635 4.030 0.960 ;
        RECT 4.200 0.950 5.085 1.120 ;
        RECT 4.200 0.425 4.370 0.950 ;
        RECT 2.505 0.255 4.370 0.425 ;
        RECT 4.540 0.085 5.080 0.780 ;
        RECT 5.755 0.085 6.085 0.640 ;
        RECT 6.755 0.085 7.085 1.130 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__o2bb2a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o2bb2ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2bb2ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.510 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.120 1.100 1.450 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.300 3.255 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.300 2.755 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.420 1.140 3.330 1.240 ;
        RECT 0.005 0.245 3.330 1.140 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.546900 ;
    PORT
      LAYER li1 ;
        RECT 1.860 1.950 2.315 2.980 ;
        RECT 1.860 1.180 2.030 1.950 ;
        RECT 1.610 1.010 2.030 1.180 ;
        RECT 1.610 0.350 1.860 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.140 1.895 0.470 3.245 ;
        RECT 0.640 1.790 0.970 2.775 ;
        RECT 1.140 1.975 1.690 3.245 ;
        RECT 2.995 1.950 3.245 3.245 ;
        RECT 0.640 1.620 1.690 1.790 ;
        RECT 1.270 1.350 1.690 1.620 ;
        RECT 1.270 0.950 1.440 1.350 ;
        RECT 0.115 0.085 0.445 0.950 ;
        RECT 0.935 0.350 1.440 0.950 ;
        RECT 2.200 0.960 3.220 1.130 ;
        RECT 2.200 0.840 2.370 0.960 ;
        RECT 2.030 0.445 2.370 0.840 ;
        RECT 2.540 0.085 2.710 0.790 ;
        RECT 2.890 0.350 3.220 0.960 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o2bb2ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2bb2ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 0.650 2.585 2.335 2.620 ;
        RECT 0.125 2.450 2.335 2.585 ;
        RECT 0.125 2.415 0.820 2.450 ;
        RECT 0.125 1.630 0.355 2.415 ;
        RECT 2.165 1.680 2.335 2.450 ;
        RECT 0.125 1.300 0.480 1.630 ;
        RECT 1.965 1.350 2.335 1.680 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 1.375 1.445 1.795 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.695 1.780 5.095 1.890 ;
        RECT 3.695 1.720 5.495 1.780 ;
        RECT 3.695 1.350 4.025 1.720 ;
        RECT 4.925 1.350 5.495 1.720 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.345 1.180 4.675 1.550 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.460 1.140 5.755 1.240 ;
        RECT 0.035 0.245 5.755 1.140 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.896000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 2.230 3.290 2.980 ;
        RECT 4.465 2.230 4.695 2.735 ;
        RECT 3.005 2.060 4.695 2.230 ;
        RECT 3.005 1.130 3.290 2.060 ;
        RECT 3.000 0.595 3.290 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 2.755 0.445 3.245 ;
        RECT 1.185 2.790 1.515 3.245 ;
        RECT 1.720 2.245 1.995 2.280 ;
        RECT 0.650 1.950 1.995 2.245 ;
        RECT 0.650 1.275 0.980 1.950 ;
        RECT 2.505 1.820 2.835 3.245 ;
        RECT 3.460 2.400 3.790 3.245 ;
        RECT 3.965 2.905 5.195 3.075 ;
        RECT 3.965 2.400 4.295 2.905 ;
        RECT 4.865 2.060 5.195 2.905 ;
        RECT 5.395 1.950 5.645 3.245 ;
        RECT 2.505 1.300 2.835 1.630 ;
        RECT 0.650 1.180 1.405 1.275 ;
        RECT 2.505 1.180 2.675 1.300 ;
        RECT 0.650 1.105 2.675 1.180 ;
        RECT 0.145 0.085 0.475 1.030 ;
        RECT 1.155 1.010 2.675 1.105 ;
        RECT 3.460 1.010 3.790 1.130 ;
        RECT 5.315 1.010 5.645 1.130 ;
        RECT 0.645 0.425 0.975 0.935 ;
        RECT 1.155 0.605 1.405 1.010 ;
        RECT 3.460 0.840 5.645 1.010 ;
        RECT 1.580 0.425 1.910 0.825 ;
        RECT 0.645 0.255 1.910 0.425 ;
        RECT 2.080 0.085 2.340 0.825 ;
        RECT 2.570 0.425 2.820 0.825 ;
        RECT 3.460 0.425 3.790 0.840 ;
        RECT 4.470 0.770 5.645 0.840 ;
        RECT 2.570 0.255 3.790 0.425 ;
        RECT 3.960 0.085 4.290 0.670 ;
        RECT 4.470 0.350 4.690 0.770 ;
        RECT 4.870 0.085 5.215 0.600 ;
        RECT 5.395 0.350 5.645 0.770 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__o2bb2ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2bb2ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.935 1.780 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.350 3.235 1.780 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.150 1.350 9.955 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.350 7.640 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 10.075 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.758400 ;
    PORT
      LAYER li1 ;
        RECT 4.155 1.970 4.485 2.980 ;
        RECT 5.055 2.150 5.305 2.980 ;
        RECT 5.055 2.120 5.635 2.150 ;
        RECT 6.495 2.120 6.825 2.735 ;
        RECT 7.395 2.120 7.725 2.735 ;
        RECT 5.055 1.970 7.725 2.120 ;
        RECT 4.155 1.950 7.725 1.970 ;
        RECT 4.155 1.800 5.715 1.950 ;
        RECT 5.545 1.130 5.715 1.800 ;
        RECT 4.695 0.960 5.885 1.130 ;
        RECT 4.695 0.595 5.025 0.960 ;
        RECT 5.545 0.595 5.885 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.105 1.950 0.355 3.245 ;
        RECT 0.555 2.120 0.885 2.980 ;
        RECT 1.085 2.290 1.255 3.245 ;
        RECT 1.455 2.120 1.785 2.980 ;
        RECT 1.985 2.290 2.155 3.245 ;
        RECT 2.355 2.120 2.685 2.980 ;
        RECT 2.885 2.290 3.055 3.245 ;
        RECT 3.255 2.120 3.585 2.980 ;
        RECT 0.555 1.950 3.585 2.120 ;
        RECT 3.415 1.630 3.585 1.950 ;
        RECT 3.785 1.820 3.955 3.245 ;
        RECT 4.685 2.140 4.855 3.245 ;
        RECT 5.505 2.320 5.835 3.245 ;
        RECT 6.045 2.905 8.110 3.075 ;
        RECT 6.045 2.290 6.310 2.905 ;
        RECT 7.010 2.290 7.210 2.905 ;
        RECT 7.910 2.120 8.110 2.905 ;
        RECT 8.295 2.290 8.560 3.245 ;
        RECT 8.745 2.120 9.075 2.980 ;
        RECT 9.260 2.290 9.465 3.245 ;
        RECT 9.645 2.120 9.975 2.980 ;
        RECT 7.910 1.950 9.975 2.120 ;
        RECT 3.415 1.300 5.375 1.630 ;
        RECT 3.415 1.180 3.605 1.300 ;
        RECT 0.115 1.010 2.095 1.180 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.055 0.350 1.235 1.010 ;
        RECT 1.415 0.085 1.745 0.840 ;
        RECT 1.925 0.425 2.095 1.010 ;
        RECT 2.275 1.010 3.605 1.180 ;
        RECT 2.275 0.595 2.605 1.010 ;
        RECT 2.775 0.425 3.105 0.840 ;
        RECT 3.275 0.595 3.605 1.010 ;
        RECT 3.785 0.425 4.035 1.130 ;
        RECT 1.925 0.255 4.035 0.425 ;
        RECT 4.265 0.425 4.515 1.130 ;
        RECT 6.065 1.010 9.965 1.180 ;
        RECT 5.205 0.425 5.375 0.790 ;
        RECT 6.065 0.425 6.235 1.010 ;
        RECT 4.265 0.255 6.235 0.425 ;
        RECT 6.415 0.085 6.745 0.830 ;
        RECT 6.915 0.350 7.165 1.010 ;
        RECT 7.345 0.085 7.675 0.830 ;
        RECT 7.845 0.350 8.095 1.010 ;
        RECT 8.275 0.085 8.605 0.830 ;
        RECT 8.785 0.350 9.035 1.010 ;
        RECT 9.205 0.085 9.535 0.830 ;
        RECT 9.715 0.350 9.965 1.010 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__o2bb2ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.300 2.775 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.445 2.275 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.445 1.435 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 0.985 1.240 ;
        RECT 0.005 0.245 2.875 1.140 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.820 0.445 2.980 ;
        RECT 0.115 0.350 0.365 1.820 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.615 2.290 1.180 3.245 ;
        RECT 1.360 2.120 1.690 2.795 ;
        RECT 0.695 1.950 1.690 2.120 ;
        RECT 2.435 1.950 2.765 3.245 ;
        RECT 0.695 1.550 0.865 1.950 ;
        RECT 0.535 1.275 0.865 1.550 ;
        RECT 0.535 1.105 1.395 1.275 ;
        RECT 0.545 0.085 0.875 0.935 ;
        RECT 1.145 0.350 1.395 1.105 ;
        RECT 1.575 0.960 2.765 1.130 ;
        RECT 1.575 0.350 1.825 0.960 ;
        RECT 2.005 0.085 2.335 0.790 ;
        RECT 2.515 0.350 2.765 0.960 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__o21a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o21a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.835 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.180 1.385 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.180 1.955 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 2.465 1.890 2.795 2.980 ;
        RECT 2.465 1.720 3.295 1.890 ;
        RECT 2.965 0.350 3.295 1.720 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.335 1.820 0.665 3.245 ;
        RECT 1.325 1.890 1.655 2.860 ;
        RECT 1.965 2.060 2.295 3.245 ;
        RECT 2.965 2.060 3.295 3.245 ;
        RECT 1.325 1.720 2.295 1.890 ;
        RECT 2.125 1.550 2.295 1.720 ;
        RECT 2.125 1.220 2.645 1.550 ;
        RECT 2.125 1.010 2.295 1.220 ;
        RECT 0.250 0.840 1.735 1.010 ;
        RECT 0.250 0.340 0.580 0.840 ;
        RECT 0.750 0.085 1.235 0.600 ;
        RECT 1.405 0.340 1.735 0.840 ;
        RECT 1.905 0.340 2.295 1.010 ;
        RECT 2.465 0.085 2.795 1.050 ;
        RECT 3.475 0.085 3.725 1.130 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o21a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.445 2.275 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.445 1.505 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.515 3.235 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 3.440 1.395 ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.890 4.145 2.980 ;
        RECT 4.815 1.890 5.145 2.980 ;
        RECT 3.815 1.780 5.145 1.890 ;
        RECT 3.815 1.720 5.635 1.780 ;
        RECT 4.965 1.550 5.635 1.720 ;
        RECT 4.965 1.005 5.135 1.550 ;
        RECT 3.990 0.835 5.135 1.005 ;
        RECT 3.990 0.330 4.240 0.835 ;
        RECT 4.965 0.350 5.135 0.835 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 1.915 0.445 3.245 ;
        RECT 0.615 2.905 1.895 3.075 ;
        RECT 0.615 1.950 0.865 2.905 ;
        RECT 1.065 2.120 1.395 2.735 ;
        RECT 1.565 2.290 1.895 2.905 ;
        RECT 2.065 2.290 2.395 3.245 ;
        RECT 2.565 2.120 2.895 2.795 ;
        RECT 3.135 2.300 3.615 3.245 ;
        RECT 1.065 1.950 3.575 2.120 ;
        RECT 4.315 2.060 4.645 3.245 ;
        RECT 5.315 1.950 5.645 3.245 ;
        RECT 3.405 1.550 3.575 1.950 ;
        RECT 3.405 1.345 4.795 1.550 ;
        RECT 0.115 1.275 0.445 1.285 ;
        RECT 0.115 1.105 2.390 1.275 ;
        RECT 0.115 0.605 0.445 1.105 ;
        RECT 0.615 0.085 0.950 0.935 ;
        RECT 1.130 0.605 1.380 1.105 ;
        RECT 1.560 0.085 1.890 0.935 ;
        RECT 2.060 0.435 2.390 1.105 ;
        RECT 2.570 1.175 4.795 1.345 ;
        RECT 2.570 0.605 2.820 1.175 ;
        RECT 3.000 0.435 3.330 1.005 ;
        RECT 2.060 0.265 3.330 0.435 ;
        RECT 3.560 0.085 3.810 1.005 ;
        RECT 4.420 0.085 4.785 0.665 ;
        RECT 5.315 0.085 5.645 1.130 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__o21a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.555 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.350 1.395 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 2.275 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.828300 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.950 1.545 2.980 ;
        RECT 0.725 1.180 0.895 1.950 ;
        RECT 0.725 1.010 2.285 1.180 ;
        RECT 1.955 0.350 2.285 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.305 1.820 0.555 3.245 ;
        RECT 1.870 1.950 2.200 3.245 ;
        RECT 0.115 0.840 0.445 1.010 ;
        RECT 0.115 0.670 1.785 0.840 ;
        RECT 0.115 0.350 0.420 0.670 ;
        RECT 0.605 0.085 1.295 0.500 ;
        RECT 1.480 0.350 1.785 0.670 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__o21ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o21ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.265 1.950 2.275 2.120 ;
        RECT 0.265 1.350 0.595 1.950 ;
        RECT 1.755 1.350 2.275 1.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.350 1.515 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.180 3.235 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.961100 ;
    PORT
      LAYER li1 ;
        RECT 1.065 2.460 1.395 2.735 ;
        RECT 2.525 2.460 2.795 2.980 ;
        RECT 1.065 2.290 2.795 2.460 ;
        RECT 2.525 1.820 2.795 2.290 ;
        RECT 2.525 1.130 2.735 1.820 ;
        RECT 2.475 0.715 2.735 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.290 0.365 3.245 ;
        RECT 0.565 2.905 1.895 3.075 ;
        RECT 0.565 2.290 0.895 2.905 ;
        RECT 1.565 2.630 1.895 2.905 ;
        RECT 2.095 2.630 2.345 3.245 ;
        RECT 2.995 1.820 3.245 3.245 ;
        RECT 0.115 1.010 2.305 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.830 ;
        RECT 1.125 0.350 1.375 1.010 ;
        RECT 1.545 0.085 1.875 0.830 ;
        RECT 2.055 0.520 2.305 1.010 ;
        RECT 2.915 0.520 3.245 1.010 ;
        RECT 2.055 0.350 3.245 0.520 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o21ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.650 1.795 1.780 ;
        RECT 0.445 1.320 1.795 1.650 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 5.635 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 3.165 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.478400 ;
    PORT
      LAYER li1 ;
        RECT 3.960 2.120 4.290 2.735 ;
        RECT 4.860 2.120 5.190 2.735 ;
        RECT 2.365 1.950 5.190 2.120 ;
        RECT 2.365 1.820 3.715 1.950 ;
        RECT 3.335 1.550 3.715 1.820 ;
        RECT 3.335 1.010 3.505 1.550 ;
        RECT 2.280 0.840 3.505 1.010 ;
        RECT 2.280 0.595 2.530 0.840 ;
        RECT 3.220 0.595 3.505 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 0.565 2.120 0.895 2.980 ;
        RECT 1.095 2.290 1.265 3.245 ;
        RECT 1.465 2.460 1.795 2.980 ;
        RECT 1.995 2.630 2.245 3.245 ;
        RECT 2.900 2.630 3.230 3.245 ;
        RECT 3.460 2.905 5.640 3.075 ;
        RECT 3.460 2.460 3.790 2.905 ;
        RECT 1.465 2.290 3.790 2.460 ;
        RECT 4.490 2.290 4.660 2.905 ;
        RECT 1.465 2.120 1.795 2.290 ;
        RECT 0.565 1.950 1.795 2.120 ;
        RECT 5.390 1.950 5.640 2.905 ;
        RECT 0.565 1.820 0.895 1.950 ;
        RECT 0.115 1.010 1.225 1.150 ;
        RECT 3.675 1.010 5.645 1.180 ;
        RECT 0.115 0.980 2.100 1.010 ;
        RECT 0.115 0.350 0.365 0.980 ;
        RECT 1.055 0.840 2.100 0.980 ;
        RECT 0.545 0.085 0.875 0.810 ;
        RECT 1.055 0.350 1.225 0.840 ;
        RECT 1.405 0.085 1.735 0.670 ;
        RECT 1.930 0.425 2.100 0.840 ;
        RECT 2.710 0.425 3.040 0.670 ;
        RECT 3.675 0.425 3.845 1.010 ;
        RECT 1.930 0.255 3.845 0.425 ;
        RECT 4.025 0.085 4.355 0.840 ;
        RECT 4.535 0.350 4.705 1.010 ;
        RECT 4.885 0.085 5.215 0.840 ;
        RECT 5.395 0.350 5.645 1.010 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__o21ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o21ba_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ba_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.130 0.550 1.800 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.130 1.315 1.800 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.180 2.845 1.550 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.065 1.140 3.830 1.240 ;
        RECT 0.005 0.245 3.830 1.140 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.820 3.755 2.980 ;
        RECT 3.585 1.130 3.755 1.820 ;
        RECT 3.390 0.350 3.755 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 1.970 0.445 3.245 ;
        RECT 1.055 2.490 1.385 2.980 ;
        RECT 1.555 2.660 1.885 3.245 ;
        RECT 2.895 2.660 3.225 3.245 ;
        RECT 1.055 2.320 3.225 2.490 ;
        RECT 1.055 1.970 1.785 2.320 ;
        RECT 1.615 1.030 1.785 1.970 ;
        RECT 1.975 1.820 2.690 2.150 ;
        RECT 1.975 1.220 2.305 1.820 ;
        RECT 3.055 1.650 3.225 2.320 ;
        RECT 3.055 1.320 3.415 1.650 ;
        RECT 0.115 0.790 1.445 0.960 ;
        RECT 0.115 0.350 0.445 0.790 ;
        RECT 0.615 0.085 0.945 0.620 ;
        RECT 1.115 0.350 1.445 0.790 ;
        RECT 1.615 0.350 1.945 1.030 ;
        RECT 2.135 1.010 2.305 1.220 ;
        RECT 2.135 0.680 2.720 1.010 ;
        RECT 2.890 0.085 3.220 1.010 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o21ba_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ba_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.180 3.735 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.720 1.180 3.235 1.550 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.505 1.050 3.835 1.240 ;
        RECT 0.005 0.245 3.835 1.050 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.010 1.820 1.440 2.070 ;
        RECT 1.010 1.130 1.180 1.820 ;
        RECT 1.010 0.350 1.340 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 2.410 0.445 2.700 ;
        RECT 0.650 2.580 0.980 3.245 ;
        RECT 1.565 2.580 2.235 3.245 ;
        RECT 2.445 2.410 2.775 2.860 ;
        RECT 0.115 2.240 2.210 2.410 ;
        RECT 0.115 1.950 0.795 2.240 ;
        RECT 0.625 1.130 0.795 1.950 ;
        RECT 1.350 1.300 1.680 1.630 ;
        RECT 1.890 1.350 2.210 2.240 ;
        RECT 2.380 1.820 2.775 2.410 ;
        RECT 3.405 1.820 3.735 3.245 ;
        RECT 0.105 0.960 0.795 1.130 ;
        RECT 1.510 1.180 1.680 1.300 ;
        RECT 2.380 1.180 2.550 1.820 ;
        RECT 1.510 1.010 2.550 1.180 ;
        RECT 0.105 0.455 0.355 0.960 ;
        RECT 0.535 0.085 0.785 0.790 ;
        RECT 1.520 0.085 1.770 0.820 ;
        RECT 1.980 0.350 2.230 1.010 ;
        RECT 3.410 0.840 3.740 1.010 ;
        RECT 2.410 0.670 3.740 0.840 ;
        RECT 2.410 0.350 2.740 0.670 ;
        RECT 2.910 0.085 3.240 0.500 ;
        RECT 3.410 0.350 3.740 0.670 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o21ba_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ba_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.175 1.450 4.675 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.845 1.450 6.115 1.780 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.180 0.835 1.550 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.925 1.240 6.235 1.395 ;
        RECT 0.035 0.245 6.235 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.093800 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.820 2.345 2.220 ;
        RECT 1.085 1.550 1.315 1.820 ;
        RECT 1.145 1.120 1.315 1.550 ;
        RECT 1.145 0.950 2.210 1.120 ;
        RECT 1.145 0.350 1.340 0.950 ;
        RECT 1.960 0.350 2.210 0.950 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.085 2.560 0.445 2.980 ;
        RECT 0.615 2.730 0.995 3.245 ;
        RECT 1.565 2.730 1.895 3.245 ;
        RECT 2.465 2.730 3.205 3.245 ;
        RECT 0.085 2.390 3.320 2.560 ;
        RECT 0.085 1.820 0.445 2.390 ;
        RECT 3.150 1.960 3.320 2.390 ;
        RECT 3.490 2.300 3.740 2.980 ;
        RECT 3.945 2.470 4.275 3.245 ;
        RECT 4.445 2.905 5.675 3.075 ;
        RECT 4.445 2.470 4.775 2.905 ;
        RECT 4.975 2.300 5.145 2.735 ;
        RECT 3.490 2.130 5.145 2.300 ;
        RECT 0.085 1.010 0.255 1.820 ;
        RECT 3.150 1.630 3.490 1.960 ;
        RECT 3.660 1.950 5.145 2.130 ;
        RECT 5.345 1.950 5.675 2.905 ;
        RECT 5.875 1.950 6.125 3.245 ;
        RECT 1.485 1.460 2.980 1.620 ;
        RECT 3.660 1.460 3.830 1.950 ;
        RECT 1.485 1.290 3.830 1.460 ;
        RECT 0.085 0.350 0.475 1.010 ;
        RECT 0.645 0.085 0.975 1.010 ;
        RECT 1.530 0.085 1.780 0.780 ;
        RECT 2.390 0.085 2.640 1.120 ;
        RECT 2.810 0.425 2.980 1.290 ;
        RECT 4.000 1.120 6.125 1.280 ;
        RECT 3.150 1.110 6.125 1.120 ;
        RECT 3.150 0.950 4.330 1.110 ;
        RECT 3.150 0.595 3.320 0.950 ;
        RECT 3.500 0.425 3.830 0.780 ;
        RECT 4.000 0.605 4.330 0.950 ;
        RECT 2.810 0.255 3.830 0.425 ;
        RECT 4.500 0.085 4.750 0.940 ;
        RECT 4.930 0.605 5.180 1.110 ;
        RECT 5.360 0.085 5.610 0.940 ;
        RECT 5.790 0.605 6.125 1.110 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__o21ba_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21bai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.300 2.775 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.630 2.275 2.890 ;
        RECT 1.750 1.300 2.275 1.630 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.565 1.780 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.980 1.050 2.875 1.240 ;
        RECT 0.005 0.245 2.875 1.050 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.475 1.990 1.840 2.980 ;
        RECT 1.305 1.820 1.840 1.990 ;
        RECT 1.305 1.130 1.475 1.820 ;
        RECT 1.085 0.350 1.475 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.135 2.120 0.465 2.980 ;
        RECT 0.635 2.290 1.305 3.245 ;
        RECT 0.135 1.950 0.915 2.120 ;
        RECT 2.520 1.950 2.770 3.245 ;
        RECT 0.745 1.630 0.915 1.950 ;
        RECT 0.745 1.300 1.135 1.630 ;
        RECT 0.745 1.280 0.915 1.300 ;
        RECT 0.110 1.110 0.915 1.280 ;
        RECT 0.110 0.350 0.360 1.110 ;
        RECT 1.645 0.960 2.765 1.130 ;
        RECT 0.540 0.085 0.870 0.940 ;
        RECT 1.645 0.350 1.815 0.960 ;
        RECT 1.995 0.085 2.335 0.680 ;
        RECT 2.515 0.350 2.765 0.960 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__o21bai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o21bai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21bai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.250 1.950 3.715 2.120 ;
        RECT 2.250 1.350 2.580 1.950 ;
        RECT 3.485 1.650 3.715 1.950 ;
        RECT 3.485 1.320 4.055 1.650 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.820 1.350 3.235 1.780 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.460 1.350 0.835 1.780 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.995 1.140 4.295 1.240 ;
        RECT 0.005 0.245 4.295 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.879200 ;
    PORT
      LAYER li1 ;
        RECT 1.530 2.460 1.780 2.980 ;
        RECT 3.050 2.460 3.220 2.735 ;
        RECT 1.530 2.290 3.220 2.460 ;
        RECT 1.530 1.180 1.865 2.290 ;
        RECT 1.615 0.615 1.865 1.180 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 1.950 0.640 2.860 ;
        RECT 0.115 1.180 0.285 1.950 ;
        RECT 1.005 1.820 1.335 3.245 ;
        RECT 1.980 2.650 2.350 3.245 ;
        RECT 2.520 2.905 3.755 3.075 ;
        RECT 2.520 2.630 2.850 2.905 ;
        RECT 3.420 2.290 3.755 2.905 ;
        RECT 3.955 1.820 4.205 3.245 ;
        RECT 1.030 1.180 1.360 1.550 ;
        RECT 0.115 1.010 1.360 1.180 ;
        RECT 2.035 1.150 3.245 1.180 ;
        RECT 2.035 1.010 4.185 1.150 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.105 0.425 1.435 0.840 ;
        RECT 2.035 0.425 2.365 1.010 ;
        RECT 3.075 0.980 4.185 1.010 ;
        RECT 1.105 0.255 2.365 0.425 ;
        RECT 2.535 0.085 2.865 0.840 ;
        RECT 3.075 0.350 3.245 0.980 ;
        RECT 3.425 0.085 3.755 0.810 ;
        RECT 3.935 0.350 4.185 0.980 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o21bai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21bai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.795 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 3.715 1.780 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.450 7.075 1.780 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.215 1.240 7.195 1.390 ;
        RECT 0.005 0.245 7.195 1.240 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.855000 ;
    PORT
      LAYER li1 ;
        RECT 2.370 2.120 2.620 2.735 ;
        RECT 3.320 2.120 3.650 2.735 ;
        RECT 4.380 2.120 4.710 2.980 ;
        RECT 2.370 2.020 4.710 2.120 ;
        RECT 5.295 2.020 5.625 2.980 ;
        RECT 2.370 1.950 5.625 2.020 ;
        RECT 3.965 1.180 4.195 1.950 ;
        RECT 4.380 1.850 5.625 1.950 ;
        RECT 3.965 1.010 5.595 1.180 ;
        RECT 4.265 0.595 4.595 1.010 ;
        RECT 5.265 0.595 5.595 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.120 2.120 0.370 2.980 ;
        RECT 0.570 2.290 0.820 3.245 ;
        RECT 1.020 2.120 1.270 2.980 ;
        RECT 1.470 2.290 1.800 3.245 ;
        RECT 2.000 2.905 4.150 3.075 ;
        RECT 2.000 2.120 2.170 2.905 ;
        RECT 2.820 2.290 3.150 2.905 ;
        RECT 3.820 2.290 4.150 2.905 ;
        RECT 4.910 2.190 5.080 3.245 ;
        RECT 5.855 2.290 6.105 3.245 ;
        RECT 6.305 2.120 6.555 2.980 ;
        RECT 0.120 1.950 2.170 2.120 ;
        RECT 2.000 1.820 2.170 1.950 ;
        RECT 5.795 1.950 6.555 2.120 ;
        RECT 6.755 2.100 7.085 3.245 ;
        RECT 5.795 1.680 5.965 1.950 ;
        RECT 4.370 1.350 5.965 1.680 ;
        RECT 5.795 1.280 5.965 1.350 ;
        RECT 0.115 1.010 3.075 1.180 ;
        RECT 5.795 1.110 6.575 1.280 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.105 0.350 1.275 1.010 ;
        RECT 1.455 0.085 1.785 0.840 ;
        RECT 1.965 0.350 2.135 1.010 ;
        RECT 2.825 0.840 3.075 1.010 ;
        RECT 2.315 0.085 2.645 0.840 ;
        RECT 2.825 0.670 4.095 0.840 ;
        RECT 2.825 0.350 3.075 0.670 ;
        RECT 3.255 0.085 3.585 0.500 ;
        RECT 3.765 0.425 4.095 0.670 ;
        RECT 4.765 0.425 5.095 0.840 ;
        RECT 5.765 0.425 6.095 0.940 ;
        RECT 6.325 0.500 6.575 1.110 ;
        RECT 3.765 0.255 6.095 0.425 ;
        RECT 6.755 0.085 7.085 1.280 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__o21bai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o22a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.235 1.470 3.715 1.800 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.470 2.995 1.800 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.335 1.470 2.005 1.800 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.585 1.305 0.670 ;
        RECT 1.085 0.255 2.470 0.585 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.400 1.420 3.210 1.465 ;
        RECT 1.400 1.410 3.800 1.420 ;
        RECT 1.400 1.240 3.835 1.410 ;
        RECT 0.005 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.675 4.030 3.520 ;
        RECT -0.190 1.660 1.160 1.675 ;
        RECT 3.190 1.660 4.030 1.675 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.445 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.365 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.615 1.985 1.850 3.245 ;
        RECT 2.395 2.140 2.725 2.980 ;
        RECT 2.175 1.970 2.725 2.140 ;
        RECT 3.385 1.970 3.715 3.245 ;
        RECT 0.425 1.300 1.095 1.630 ;
        RECT 2.175 1.300 2.345 1.970 ;
        RECT 0.925 1.130 2.345 1.300 ;
        RECT 1.905 1.105 2.345 1.130 ;
        RECT 2.535 1.130 3.725 1.300 ;
        RECT 0.545 0.085 0.875 0.960 ;
        RECT 2.535 0.935 2.705 1.130 ;
        RECT 1.475 0.755 2.705 0.935 ;
        RECT 2.885 0.085 3.225 0.960 ;
        RECT 3.395 0.630 3.725 1.130 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o22a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o22a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o22a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.300 3.735 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.710 1.430 3.235 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.430 1.875 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.430 2.500 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.820 0.965 2.980 ;
        RECT 0.635 1.130 0.805 1.820 ;
        RECT 0.535 0.820 0.865 1.130 ;
        RECT 0.535 0.350 0.790 0.820 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.135 1.820 0.465 3.245 ;
        RECT 1.135 2.290 1.790 3.245 ;
        RECT 2.350 2.120 2.680 2.940 ;
        RECT 1.135 1.950 2.680 2.120 ;
        RECT 3.400 1.950 3.730 3.245 ;
        RECT 1.135 1.630 1.305 1.950 ;
        RECT 0.975 1.300 1.305 1.630 ;
        RECT 1.135 1.130 1.305 1.300 ;
        RECT 0.105 0.085 0.365 1.130 ;
        RECT 1.135 0.880 2.295 1.130 ;
        RECT 2.005 0.800 2.295 0.880 ;
        RECT 2.465 0.960 3.725 1.130 ;
        RECT 0.965 0.085 1.295 0.640 ;
        RECT 1.505 0.520 1.835 0.710 ;
        RECT 2.465 0.520 2.795 0.960 ;
        RECT 1.505 0.350 2.795 0.520 ;
        RECT 2.965 0.085 3.295 0.790 ;
        RECT 3.475 0.350 3.725 0.960 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o22a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o22a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o22a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.450 2.275 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.450 1.515 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.570 2.275 0.670 ;
        RECT 2.045 0.255 2.610 0.570 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.450 3.505 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 4.350 1.450 ;
        RECT 0.005 0.245 6.715 1.240 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.125600 ;
    PORT
      LAYER li1 ;
        RECT 4.600 2.020 4.930 2.980 ;
        RECT 5.775 2.020 6.105 2.980 ;
        RECT 4.600 1.850 6.105 2.020 ;
        RECT 5.935 1.410 6.105 1.850 ;
        RECT 5.935 1.180 6.595 1.410 ;
        RECT 4.980 1.010 6.105 1.180 ;
        RECT 4.980 0.350 5.230 1.010 ;
        RECT 5.920 0.350 6.105 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.115 1.940 0.365 3.245 ;
        RECT 0.565 2.905 1.895 3.075 ;
        RECT 0.565 1.950 0.895 2.905 ;
        RECT 1.065 2.120 1.395 2.735 ;
        RECT 1.565 2.290 1.895 2.905 ;
        RECT 2.065 2.290 2.395 3.245 ;
        RECT 2.565 2.905 3.895 3.075 ;
        RECT 2.565 2.290 2.895 2.905 ;
        RECT 3.065 2.120 3.395 2.735 ;
        RECT 3.565 2.290 3.895 2.905 ;
        RECT 1.065 1.950 3.845 2.120 ;
        RECT 3.675 1.680 3.845 1.950 ;
        RECT 4.100 1.850 4.430 3.245 ;
        RECT 5.200 2.190 5.530 3.245 ;
        RECT 6.275 1.820 6.605 3.245 ;
        RECT 3.675 1.510 5.765 1.680 ;
        RECT 4.415 1.350 5.765 1.510 ;
        RECT 0.115 1.280 0.445 1.340 ;
        RECT 3.910 1.280 4.240 1.340 ;
        RECT 0.115 1.110 4.240 1.280 ;
        RECT 0.115 0.660 0.445 1.110 ;
        RECT 0.615 0.085 0.945 0.940 ;
        RECT 1.125 0.660 1.375 1.110 ;
        RECT 2.045 1.090 4.240 1.110 ;
        RECT 1.545 0.085 1.875 0.940 ;
        RECT 2.045 0.840 2.375 1.090 ;
        RECT 4.415 0.920 4.585 1.350 ;
        RECT 2.545 0.750 4.585 0.920 ;
        RECT 2.545 0.740 3.810 0.750 ;
        RECT 3.480 0.660 3.810 0.740 ;
        RECT 4.470 0.085 4.800 0.580 ;
        RECT 5.410 0.085 5.740 0.790 ;
        RECT 6.275 0.085 6.605 1.010 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__o22a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o22ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.300 2.775 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.350 1.865 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.180 0.445 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.350 1.315 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.780 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.895900 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.950 1.550 2.980 ;
        RECT 0.625 1.130 0.795 1.950 ;
        RECT 0.615 0.655 1.065 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.125 1.820 0.455 3.245 ;
        RECT 2.255 1.950 2.585 3.245 ;
        RECT 0.115 0.485 0.445 1.010 ;
        RECT 1.340 0.960 2.670 1.130 ;
        RECT 1.340 0.485 1.670 0.960 ;
        RECT 0.115 0.315 1.670 0.485 ;
        RECT 1.840 0.085 2.170 0.790 ;
        RECT 2.340 0.350 2.670 0.960 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__o22ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o22ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o22ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.910 1.350 4.675 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.630 3.715 1.780 ;
        RECT 2.665 1.390 3.715 1.630 ;
        RECT 2.665 1.300 3.335 1.390 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.315 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.350 1.815 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.212200 ;
    PORT
      LAYER li1 ;
        RECT 1.570 2.120 1.800 2.735 ;
        RECT 1.570 1.970 2.275 2.120 ;
        RECT 3.060 1.970 3.310 2.735 ;
        RECT 1.570 1.950 3.310 1.970 ;
        RECT 2.045 1.800 3.310 1.950 ;
        RECT 2.045 1.180 2.275 1.800 ;
        RECT 0.615 1.010 2.275 1.180 ;
        RECT 0.615 0.595 0.945 1.010 ;
        RECT 1.615 0.595 1.945 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.120 2.120 0.370 2.980 ;
        RECT 0.570 2.290 0.900 3.245 ;
        RECT 1.070 2.905 2.300 3.075 ;
        RECT 1.070 2.120 1.400 2.905 ;
        RECT 1.970 2.290 2.300 2.905 ;
        RECT 2.530 2.905 3.680 3.075 ;
        RECT 2.530 2.140 2.860 2.905 ;
        RECT 0.120 1.950 1.400 2.120 ;
        RECT 3.510 2.120 3.680 2.905 ;
        RECT 3.880 2.290 4.130 3.245 ;
        RECT 4.330 2.120 4.660 2.980 ;
        RECT 3.510 1.950 4.660 2.120 ;
        RECT 3.505 1.130 4.685 1.180 ;
        RECT 0.115 0.425 0.445 1.130 ;
        RECT 2.455 1.010 4.685 1.130 ;
        RECT 2.455 0.960 3.755 1.010 ;
        RECT 2.455 0.840 2.785 0.960 ;
        RECT 1.115 0.425 1.445 0.840 ;
        RECT 2.115 0.425 2.785 0.840 ;
        RECT 0.115 0.255 2.785 0.425 ;
        RECT 2.955 0.085 3.285 0.790 ;
        RECT 3.505 0.350 3.755 0.960 ;
        RECT 3.925 0.085 4.255 0.840 ;
        RECT 4.435 0.350 4.685 1.010 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o22ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o22ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.890 3.235 2.150 ;
        RECT 1.380 1.720 3.810 1.890 ;
        RECT 1.380 1.650 1.550 1.720 ;
        RECT 0.540 1.320 1.550 1.650 ;
        RECT 3.640 1.680 3.810 1.720 ;
        RECT 3.640 1.350 3.970 1.680 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.180 3.235 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.290 1.300 5.635 1.630 ;
        RECT 5.405 1.260 5.635 1.300 ;
        RECT 7.400 1.260 7.730 1.550 ;
        RECT 5.405 1.090 7.730 1.260 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.680 7.155 1.780 ;
        RECT 5.805 1.430 7.155 1.680 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 8.155 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.388000 ;
    PORT
      LAYER li1 ;
        RECT 2.020 2.320 4.150 2.490 ;
        RECT 2.020 2.060 2.350 2.320 ;
        RECT 3.980 2.020 4.150 2.320 ;
        RECT 5.770 2.120 6.100 2.735 ;
        RECT 6.670 2.120 7.000 2.735 ;
        RECT 5.770 2.020 8.070 2.120 ;
        RECT 3.980 1.950 8.070 2.020 ;
        RECT 3.980 1.850 6.100 1.950 ;
        RECT 4.405 0.920 5.155 1.130 ;
        RECT 7.900 0.920 8.070 1.950 ;
        RECT 4.405 0.750 8.070 0.920 ;
        RECT 6.205 0.595 6.535 0.750 ;
        RECT 7.205 0.595 7.535 0.750 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.120 1.820 0.370 3.245 ;
        RECT 0.570 2.230 0.850 2.980 ;
        RECT 1.020 2.400 1.350 3.245 ;
        RECT 1.520 2.660 3.700 2.980 ;
        RECT 3.870 2.660 4.200 3.245 ;
        RECT 1.520 2.230 1.850 2.660 ;
        RECT 0.570 2.060 1.850 2.230 ;
        RECT 4.370 2.360 4.700 2.980 ;
        RECT 4.900 2.530 5.150 3.245 ;
        RECT 5.320 2.905 7.500 3.075 ;
        RECT 5.320 2.360 5.570 2.905 ;
        RECT 4.370 2.190 5.570 2.360 ;
        RECT 6.300 2.290 6.470 2.905 ;
        RECT 7.170 2.290 7.500 2.905 ;
        RECT 7.670 2.290 8.000 3.245 ;
        RECT 0.570 1.820 0.900 2.060 ;
        RECT 0.115 1.010 1.375 1.150 ;
        RECT 3.905 1.010 4.235 1.130 ;
        RECT 0.115 0.980 4.235 1.010 ;
        RECT 0.115 0.350 0.445 0.980 ;
        RECT 1.125 0.840 4.235 0.980 ;
        RECT 0.615 0.085 0.945 0.810 ;
        RECT 1.125 0.350 1.375 0.840 ;
        RECT 1.545 0.085 1.875 0.670 ;
        RECT 2.055 0.350 2.305 0.840 ;
        RECT 2.475 0.085 2.805 0.670 ;
        RECT 2.985 0.350 3.235 0.840 ;
        RECT 3.405 0.085 3.735 0.670 ;
        RECT 3.905 0.580 4.235 0.840 ;
        RECT 3.905 0.425 6.035 0.580 ;
        RECT 6.705 0.425 7.035 0.580 ;
        RECT 7.715 0.425 8.045 0.580 ;
        RECT 3.905 0.255 8.045 0.425 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__o22ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o31a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o31a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.350 1.315 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.300 1.835 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.375 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.350 2.915 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.455 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.445 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.625 2.290 1.090 3.245 ;
        RECT 2.195 2.120 2.525 2.880 ;
        RECT 2.735 2.290 3.050 3.245 ;
        RECT 0.625 1.950 3.255 2.120 ;
        RECT 0.625 1.650 0.795 1.950 ;
        RECT 0.425 1.320 0.795 1.650 ;
        RECT 3.085 1.130 3.255 1.950 ;
        RECT 0.615 0.085 0.945 1.130 ;
        RECT 1.125 0.960 2.745 1.130 ;
        RECT 1.125 0.450 1.460 0.960 ;
        RECT 1.765 0.085 2.130 0.780 ;
        RECT 2.415 0.450 2.745 0.960 ;
        RECT 2.915 0.450 3.255 1.130 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o31a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o31a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o31a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.350 1.795 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.470 2.315 2.150 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.180 2.885 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.300 3.725 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.604800 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.820 0.950 2.150 ;
        RECT 0.775 1.130 0.945 1.820 ;
        RECT 0.615 0.350 0.945 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 2.660 0.445 3.245 ;
        RECT 1.070 2.660 1.595 3.245 ;
        RECT 2.765 2.490 3.225 2.980 ;
        RECT 0.225 2.320 3.225 2.490 ;
        RECT 0.225 1.650 0.395 2.320 ;
        RECT 2.765 1.940 3.225 2.320 ;
        RECT 3.395 1.950 3.725 3.245 ;
        RECT 0.225 1.320 0.605 1.650 ;
        RECT 3.055 1.130 3.225 1.940 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 1.115 0.085 1.445 1.130 ;
        RECT 1.615 0.940 1.945 1.130 ;
        RECT 3.055 0.960 3.725 1.130 ;
        RECT 1.615 0.790 2.850 0.940 ;
        RECT 1.615 0.770 3.225 0.790 ;
        RECT 1.615 0.350 1.945 0.770 ;
        RECT 2.115 0.085 2.510 0.600 ;
        RECT 2.680 0.460 3.225 0.770 ;
        RECT 3.395 0.350 3.725 0.960 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o31a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o31a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o31a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.455 5.875 1.785 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.115 1.455 6.595 1.785 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.455 5.155 1.785 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.470 3.235 2.150 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.330 1.240 6.690 1.395 ;
        RECT 0.035 0.245 6.690 1.240 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.970 0.835 2.980 ;
        RECT 1.480 1.970 1.810 2.980 ;
        RECT 0.575 1.800 1.810 1.970 ;
        RECT 0.575 1.130 0.835 1.800 ;
        RECT 0.575 0.960 1.700 1.130 ;
        RECT 0.575 0.350 0.905 0.960 ;
        RECT 1.450 0.350 1.700 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.130 1.820 0.380 3.245 ;
        RECT 1.030 2.140 1.280 3.245 ;
        RECT 2.010 1.820 2.260 3.245 ;
        RECT 2.465 2.545 2.715 2.980 ;
        RECT 2.915 2.715 3.245 3.245 ;
        RECT 3.925 2.545 4.255 2.980 ;
        RECT 2.465 2.375 4.255 2.545 ;
        RECT 2.465 1.630 2.715 2.375 ;
        RECT 4.435 2.205 4.645 2.980 ;
        RECT 4.825 2.465 5.075 2.980 ;
        RECT 5.275 2.635 5.605 3.245 ;
        RECT 5.775 2.465 6.105 2.980 ;
        RECT 4.825 2.295 6.105 2.465 ;
        RECT 3.475 2.125 4.645 2.205 ;
        RECT 6.275 2.125 6.605 2.980 ;
        RECT 3.475 1.955 6.605 2.125 ;
        RECT 1.005 1.300 2.715 1.630 ;
        RECT 2.545 1.130 3.270 1.300 ;
        RECT 0.145 0.085 0.395 1.130 ;
        RECT 1.085 0.085 1.255 0.790 ;
        RECT 1.880 0.085 2.210 1.130 ;
        RECT 2.440 0.435 2.770 0.960 ;
        RECT 2.940 0.605 3.270 1.130 ;
        RECT 3.450 1.115 6.580 1.285 ;
        RECT 3.450 0.435 3.780 1.115 ;
        RECT 2.440 0.265 3.780 0.435 ;
        RECT 3.960 0.085 4.210 0.945 ;
        RECT 4.390 0.605 4.640 1.115 ;
        RECT 4.820 0.085 5.150 0.945 ;
        RECT 5.320 0.605 5.570 1.115 ;
        RECT 5.750 0.085 6.080 0.945 ;
        RECT 6.250 0.605 6.580 1.115 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__o31a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o31ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o31ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.300 1.180 2.890 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.690 1.350 2.275 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.300 2.775 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.875 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.020700 ;
    PORT
      LAYER li1 ;
        RECT 1.350 1.950 2.230 2.980 ;
        RECT 1.350 1.130 1.520 1.950 ;
        RECT 1.350 0.960 2.765 1.130 ;
        RECT 2.435 0.350 2.765 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.130 1.820 0.380 3.245 ;
        RECT 2.410 1.950 2.740 3.245 ;
        RECT 0.115 0.085 0.445 1.010 ;
        RECT 0.625 0.790 0.875 1.130 ;
        RECT 0.625 0.620 2.265 0.790 ;
        RECT 0.625 0.350 0.875 0.620 ;
        RECT 1.055 0.085 1.755 0.450 ;
        RECT 1.935 0.350 2.265 0.620 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__o31ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o31ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o31ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.315 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 2.275 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 3.445 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.685 1.350 4.695 1.680 ;
        RECT 4.365 1.180 4.695 1.350 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.790 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.297000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 2.120 2.755 2.735 ;
        RECT 3.455 2.120 3.785 2.980 ;
        RECT 2.505 2.020 3.785 2.120 ;
        RECT 4.355 2.020 4.685 2.980 ;
        RECT 2.505 1.950 4.685 2.020 ;
        RECT 2.505 1.820 2.835 1.950 ;
        RECT 3.615 1.850 4.685 1.950 ;
        RECT 2.665 1.180 2.835 1.820 ;
        RECT 2.665 1.010 4.180 1.180 ;
        RECT 3.850 0.610 4.180 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.120 2.120 0.370 2.980 ;
        RECT 0.570 2.290 0.820 3.245 ;
        RECT 1.020 2.120 1.350 2.980 ;
        RECT 1.550 2.905 3.285 3.075 ;
        RECT 1.550 2.290 1.720 2.905 ;
        RECT 1.920 2.120 2.250 2.735 ;
        RECT 2.955 2.290 3.285 2.905 ;
        RECT 3.985 2.190 4.155 3.245 ;
        RECT 0.120 1.950 2.250 2.120 ;
        RECT 0.115 1.010 2.445 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.825 ;
        RECT 1.115 0.350 1.445 1.010 ;
        RECT 2.115 0.840 2.445 1.010 ;
        RECT 1.615 0.085 1.945 0.825 ;
        RECT 2.115 0.670 3.670 0.840 ;
        RECT 2.115 0.350 2.445 0.670 ;
        RECT 2.625 0.085 3.240 0.500 ;
        RECT 3.420 0.425 3.670 0.670 ;
        RECT 4.350 0.425 4.680 1.010 ;
        RECT 3.420 0.255 4.680 0.425 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o31ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o31ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.795 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 3.715 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.835 1.350 6.115 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.350 7.790 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 8.635 1.280 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.803200 ;
    PORT
      LAYER li1 ;
        RECT 4.700 2.150 4.970 2.735 ;
        RECT 3.965 2.120 4.970 2.150 ;
        RECT 5.600 2.120 5.930 2.735 ;
        RECT 6.550 2.120 6.880 2.980 ;
        RECT 8.195 2.120 8.525 2.980 ;
        RECT 3.965 1.950 8.525 2.120 ;
        RECT 3.965 1.550 4.665 1.950 ;
        RECT 8.195 1.820 8.525 1.950 ;
        RECT 4.495 1.180 4.665 1.550 ;
        RECT 4.495 1.010 8.095 1.180 ;
        RECT 6.905 0.920 8.095 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.120 2.120 0.370 2.980 ;
        RECT 0.570 2.290 0.900 3.245 ;
        RECT 1.100 2.120 1.270 2.980 ;
        RECT 1.470 2.290 1.800 3.245 ;
        RECT 1.970 2.120 2.300 2.980 ;
        RECT 2.470 2.905 6.380 3.075 ;
        RECT 2.470 2.290 2.800 2.905 ;
        RECT 2.970 2.540 3.300 2.735 ;
        RECT 3.640 2.710 3.970 2.905 ;
        RECT 4.140 2.540 4.470 2.735 ;
        RECT 2.970 2.370 4.470 2.540 ;
        RECT 2.970 2.120 3.300 2.370 ;
        RECT 5.150 2.290 5.400 2.905 ;
        RECT 6.130 2.290 6.380 2.905 ;
        RECT 7.050 2.290 8.025 3.245 ;
        RECT 0.120 1.950 3.300 2.120 ;
        RECT 1.970 1.820 2.300 1.950 ;
        RECT 0.115 1.010 4.325 1.180 ;
        RECT 0.115 0.920 2.305 1.010 ;
        RECT 0.115 0.390 0.445 0.920 ;
        RECT 0.615 0.085 0.945 0.750 ;
        RECT 1.475 0.085 1.805 0.750 ;
        RECT 1.975 0.390 2.305 0.920 ;
        RECT 2.495 0.085 2.960 0.805 ;
        RECT 3.145 0.390 3.475 1.010 ;
        RECT 4.155 0.840 4.325 1.010 ;
        RECT 3.645 0.085 3.975 0.840 ;
        RECT 4.155 0.750 5.775 0.840 ;
        RECT 4.155 0.670 6.805 0.750 ;
        RECT 4.155 0.390 4.325 0.670 ;
        RECT 5.445 0.580 6.805 0.670 ;
        RECT 4.585 0.085 5.265 0.500 ;
        RECT 5.445 0.390 5.775 0.580 ;
        RECT 6.475 0.560 6.805 0.580 ;
        RECT 7.335 0.560 7.665 0.750 ;
        RECT 8.265 0.560 8.525 1.170 ;
        RECT 5.955 0.085 6.295 0.410 ;
        RECT 6.475 0.390 8.525 0.560 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__o31ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o32a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o32a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.350 1.315 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.350 1.825 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.350 2.365 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.410 1.180 3.735 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.535 1.350 2.895 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 1.140 1.065 1.240 ;
        RECT 0.120 0.245 3.815 1.140 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.445 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.560 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.615 2.290 0.945 3.245 ;
        RECT 2.205 2.120 2.595 2.880 ;
        RECT 3.320 2.290 3.650 3.245 ;
        RECT 0.615 1.950 3.235 2.120 ;
        RECT 3.410 1.970 3.650 2.290 ;
        RECT 0.615 1.650 0.785 1.950 ;
        RECT 0.425 1.320 0.785 1.650 ;
        RECT 3.065 1.180 3.235 1.950 ;
        RECT 0.730 0.085 1.060 1.030 ;
        RECT 1.230 1.010 2.560 1.180 ;
        RECT 1.230 0.350 1.560 1.010 ;
        RECT 1.730 0.085 2.060 0.820 ;
        RECT 2.230 0.520 2.560 1.010 ;
        RECT 2.730 1.010 3.235 1.180 ;
        RECT 2.730 0.700 3.225 1.010 ;
        RECT 3.405 0.520 3.655 1.010 ;
        RECT 2.230 0.340 3.655 0.520 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o32a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o32a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o32a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.350 1.795 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.350 2.315 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 2.855 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 4.355 1.180 4.685 2.890 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.350 3.715 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.820 0.895 2.980 ;
        RECT 0.535 1.130 0.705 1.820 ;
        RECT 0.535 0.960 1.050 1.130 ;
        RECT 0.720 0.350 1.050 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.065 2.290 1.600 3.245 ;
        RECT 2.675 2.120 3.110 2.880 ;
        RECT 3.815 2.290 4.145 3.245 ;
        RECT 1.065 1.950 4.185 2.120 ;
        RECT 1.065 1.650 1.235 1.950 ;
        RECT 0.875 1.320 1.235 1.650 ;
        RECT 0.115 0.790 0.365 1.140 ;
        RECT 0.115 0.085 0.540 0.790 ;
        RECT 1.220 0.085 1.550 1.130 ;
        RECT 1.720 1.010 3.050 1.180 ;
        RECT 4.015 1.045 4.185 1.950 ;
        RECT 1.720 0.350 2.050 1.010 ;
        RECT 2.220 0.085 2.550 0.840 ;
        RECT 2.720 0.520 3.050 1.010 ;
        RECT 3.220 0.715 4.185 1.045 ;
        RECT 4.355 0.520 4.615 1.010 ;
        RECT 2.720 0.350 4.615 0.520 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o32a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o32a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o32a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.120 7.295 1.410 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.075 1.780 6.405 1.800 ;
        RECT 6.075 1.580 8.035 1.780 ;
        RECT 6.075 1.130 6.405 1.580 ;
        RECT 7.565 1.450 8.035 1.580 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.065 1.180 5.735 1.510 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.685 2.360 5.905 2.530 ;
        RECT 2.685 1.780 2.855 2.360 ;
        RECT 5.735 1.850 5.905 2.360 ;
        RECT 2.525 1.450 2.855 1.780 ;
        RECT 4.495 1.680 5.905 1.850 ;
        RECT 4.495 1.450 4.825 1.680 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.925 1.270 4.255 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.180 1.160 2.680 1.240 ;
        RECT 0.075 1.140 2.680 1.160 ;
        RECT 0.075 0.245 8.155 1.140 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.313300 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.950 0.895 2.980 ;
        RECT 1.565 1.950 1.895 2.980 ;
        RECT 0.565 1.780 1.895 1.950 ;
        RECT 0.565 1.650 0.895 1.780 ;
        RECT 0.125 1.480 0.895 1.650 ;
        RECT 0.125 1.310 0.355 1.480 ;
        RECT 0.125 1.140 1.015 1.310 ;
        RECT 0.685 1.110 1.015 1.140 ;
        RECT 0.685 0.940 2.015 1.110 ;
        RECT 0.685 0.350 1.015 0.940 ;
        RECT 1.685 0.350 2.015 0.940 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.065 2.120 1.395 3.245 ;
        RECT 2.085 1.950 2.415 3.245 ;
        RECT 2.655 2.700 4.025 2.960 ;
        RECT 4.195 2.700 4.525 3.245 ;
        RECT 4.785 2.700 6.245 2.980 ;
        RECT 6.805 2.730 7.135 3.245 ;
        RECT 6.075 2.560 6.245 2.700 ;
        RECT 7.715 2.560 8.045 2.980 ;
        RECT 6.075 2.390 8.045 2.560 ;
        RECT 6.155 2.200 6.675 2.220 ;
        RECT 3.230 2.020 5.565 2.190 ;
        RECT 3.230 1.920 3.575 2.020 ;
        RECT 6.155 1.970 7.595 2.200 ;
        RECT 7.265 1.950 7.595 1.970 ;
        RECT 7.765 1.950 8.045 2.390 ;
        RECT 1.255 1.280 2.355 1.610 ;
        RECT 3.230 1.280 3.560 1.920 ;
        RECT 2.185 1.110 3.560 1.280 ;
        RECT 3.300 1.100 3.560 1.110 ;
        RECT 0.185 0.085 0.515 0.970 ;
        RECT 1.185 0.085 1.515 0.770 ;
        RECT 2.240 0.085 2.570 0.940 ;
        RECT 2.800 0.425 3.130 0.940 ;
        RECT 3.300 0.930 4.560 1.100 ;
        RECT 3.300 0.595 3.560 0.930 ;
        RECT 3.730 0.425 4.060 0.760 ;
        RECT 4.230 0.595 4.560 0.930 ;
        RECT 4.730 0.960 5.060 1.010 ;
        RECT 4.730 0.950 6.060 0.960 ;
        RECT 7.715 0.950 8.045 1.030 ;
        RECT 4.730 0.790 8.045 0.950 ;
        RECT 4.730 0.425 5.060 0.790 ;
        RECT 5.730 0.780 8.045 0.790 ;
        RECT 2.800 0.255 5.060 0.425 ;
        RECT 5.230 0.085 5.560 0.620 ;
        RECT 5.730 0.350 6.060 0.780 ;
        RECT 6.230 0.085 6.560 0.610 ;
        RECT 6.740 0.350 6.990 0.780 ;
        RECT 7.160 0.085 7.545 0.600 ;
        RECT 7.715 0.350 8.045 0.780 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__o32a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o32ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o32ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.880 1.180 3.235 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.445 2.890 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 2.520 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.180 0.445 1.550 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.350 1.315 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.250 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.992900 ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.950 1.375 2.980 ;
        RECT 0.635 1.130 0.805 1.950 ;
        RECT 0.615 0.720 1.140 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.135 1.820 0.465 3.245 ;
        RECT 2.835 1.820 3.165 3.245 ;
        RECT 1.350 1.010 2.710 1.180 ;
        RECT 0.115 0.520 0.445 1.010 ;
        RECT 1.350 0.520 1.680 1.010 ;
        RECT 0.115 0.350 1.680 0.520 ;
        RECT 1.850 0.085 2.180 0.810 ;
        RECT 2.380 0.350 2.710 1.010 ;
        RECT 2.880 0.085 3.140 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o32ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o32ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.195 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.755 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.350 1.815 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.315 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 6.235 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.138200 ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.120 0.895 2.735 ;
        RECT 2.925 2.120 3.255 2.735 ;
        RECT 0.565 1.950 3.255 2.120 ;
        RECT 2.925 1.820 3.255 1.950 ;
        RECT 2.925 1.180 3.095 1.820 ;
        RECT 0.545 1.010 3.095 1.180 ;
        RECT 0.545 0.610 0.875 1.010 ;
        RECT 1.545 0.610 1.875 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.115 2.905 1.265 3.075 ;
        RECT 0.115 1.950 0.365 2.905 ;
        RECT 1.095 2.460 1.265 2.905 ;
        RECT 1.465 2.630 1.715 3.245 ;
        RECT 1.915 2.460 2.245 2.980 ;
        RECT 1.095 2.290 2.245 2.460 ;
        RECT 2.475 2.905 4.605 3.075 ;
        RECT 2.475 2.290 2.725 2.905 ;
        RECT 3.455 1.950 3.625 2.905 ;
        RECT 3.825 2.120 4.075 2.735 ;
        RECT 4.275 2.290 4.605 2.905 ;
        RECT 4.835 2.290 5.165 3.245 ;
        RECT 5.335 2.120 5.670 2.980 ;
        RECT 3.825 1.950 5.670 2.120 ;
        RECT 5.870 1.950 6.120 3.245 ;
        RECT 0.115 0.425 0.365 1.130 ;
        RECT 3.305 1.010 6.125 1.180 ;
        RECT 3.305 0.840 3.635 1.010 ;
        RECT 1.045 0.425 1.375 0.825 ;
        RECT 2.045 0.670 3.635 0.840 ;
        RECT 2.045 0.425 2.375 0.670 ;
        RECT 0.115 0.255 2.375 0.425 ;
        RECT 2.555 0.085 3.125 0.500 ;
        RECT 3.305 0.350 3.635 0.670 ;
        RECT 3.805 0.085 4.135 0.800 ;
        RECT 4.305 0.350 4.635 1.010 ;
        RECT 4.805 0.085 5.625 0.805 ;
        RECT 5.795 0.350 6.125 1.010 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__o32ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o32ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.350 10.915 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.350 8.515 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.430 5.635 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.430 4.195 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.430 1.795 1.780 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 10.780 1.240 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.287500 ;
    PORT
      LAYER li1 ;
        RECT 0.645 2.120 0.815 2.735 ;
        RECT 1.465 2.120 1.795 2.735 ;
        RECT 4.735 2.120 5.065 2.735 ;
        RECT 5.635 2.120 5.965 2.735 ;
        RECT 0.645 1.950 5.975 2.120 ;
        RECT 5.805 1.260 5.975 1.950 ;
        RECT 0.545 1.090 5.975 1.260 ;
        RECT 0.545 0.595 0.875 1.090 ;
        RECT 1.555 0.595 1.805 1.090 ;
        RECT 2.475 0.595 2.805 1.090 ;
        RECT 3.475 0.595 3.805 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.115 2.905 2.245 3.075 ;
        RECT 0.115 1.950 0.445 2.905 ;
        RECT 1.015 2.290 1.265 2.905 ;
        RECT 1.995 2.460 2.245 2.905 ;
        RECT 2.445 2.630 2.615 3.245 ;
        RECT 2.815 2.460 3.145 2.980 ;
        RECT 3.345 2.630 3.515 3.245 ;
        RECT 3.725 2.460 4.055 2.980 ;
        RECT 1.995 2.290 4.055 2.460 ;
        RECT 4.285 2.905 8.465 3.075 ;
        RECT 4.285 2.290 4.535 2.905 ;
        RECT 5.265 2.290 5.435 2.905 ;
        RECT 6.145 1.950 6.465 2.905 ;
        RECT 6.635 2.120 6.965 2.735 ;
        RECT 7.135 2.290 7.465 2.905 ;
        RECT 7.635 2.120 7.965 2.735 ;
        RECT 8.135 2.290 8.465 2.905 ;
        RECT 8.695 2.290 8.945 3.245 ;
        RECT 9.145 2.120 9.475 2.980 ;
        RECT 9.645 2.290 9.975 3.245 ;
        RECT 10.145 2.120 10.475 2.980 ;
        RECT 6.635 1.950 10.475 2.120 ;
        RECT 10.675 1.950 10.925 3.245 ;
        RECT 0.115 0.425 0.365 1.130 ;
        RECT 6.330 1.010 10.670 1.180 ;
        RECT 6.330 0.920 6.670 1.010 ;
        RECT 1.045 0.425 1.375 0.920 ;
        RECT 1.975 0.425 2.305 0.920 ;
        RECT 2.975 0.425 3.305 0.920 ;
        RECT 3.975 0.750 6.670 0.920 ;
        RECT 3.975 0.425 4.305 0.750 ;
        RECT 0.115 0.255 4.305 0.425 ;
        RECT 4.485 0.085 4.815 0.580 ;
        RECT 4.995 0.330 5.325 0.750 ;
        RECT 5.495 0.085 5.825 0.580 ;
        RECT 5.995 0.330 6.670 0.750 ;
        RECT 6.840 0.085 7.170 0.840 ;
        RECT 7.340 0.350 7.670 1.010 ;
        RECT 7.840 0.085 8.170 0.840 ;
        RECT 8.340 0.350 8.670 1.010 ;
        RECT 8.840 0.085 9.170 0.840 ;
        RECT 9.340 0.350 9.670 1.010 ;
        RECT 9.840 0.085 10.170 0.840 ;
        RECT 10.340 0.350 10.670 1.010 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__o32ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o41a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o41a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 3.610 1.350 4.195 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.300 3.370 2.890 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 2.470 1.220 2.800 2.890 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.264000 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.190 2.275 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.450 1.580 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 1.055 1.240 ;
        RECT 0.005 0.245 4.315 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.290 0.445 2.980 ;
        RECT 0.115 1.130 0.285 2.290 ;
        RECT 0.115 0.350 0.375 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.615 2.290 1.540 3.245 ;
        RECT 1.750 2.120 2.080 2.845 ;
        RECT 3.760 2.320 4.205 3.245 ;
        RECT 0.455 1.950 2.080 2.120 ;
        RECT 0.455 1.350 0.785 1.950 ;
        RECT 0.615 1.280 0.785 1.350 ;
        RECT 0.615 1.110 1.505 1.280 ;
        RECT 0.545 0.085 0.945 0.940 ;
        RECT 1.175 0.350 1.505 1.110 ;
        RECT 3.875 1.020 4.205 1.030 ;
        RECT 1.675 0.850 4.205 1.020 ;
        RECT 1.675 0.350 2.005 0.850 ;
        RECT 2.175 0.085 2.505 0.680 ;
        RECT 2.675 0.350 3.005 0.850 ;
        RECT 3.175 0.085 3.705 0.680 ;
        RECT 3.875 0.350 4.205 0.850 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o41a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o41a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o41a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.595 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.920 1.315 2.890 ;
        RECT 0.835 1.350 1.165 1.920 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.680 1.795 2.890 ;
        RECT 1.405 1.350 1.795 1.680 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.350 2.305 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 3.235 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.950 1.410 4.155 2.980 ;
        RECT 3.950 1.180 4.195 1.410 ;
        RECT 3.950 1.130 4.185 1.180 ;
        RECT 3.855 0.350 4.185 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 1.950 0.445 3.245 ;
        RECT 2.125 2.120 2.455 2.980 ;
        RECT 2.695 2.290 3.780 3.245 ;
        RECT 2.125 1.950 3.735 2.120 ;
        RECT 3.405 1.300 3.735 1.950 ;
        RECT 4.355 1.820 4.685 3.245 ;
        RECT 3.405 1.180 3.575 1.300 ;
        RECT 0.115 1.010 2.625 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.115 0.350 1.445 1.010 ;
        RECT 1.615 0.085 2.125 0.815 ;
        RECT 2.295 0.350 2.625 1.010 ;
        RECT 2.795 1.010 3.575 1.180 ;
        RECT 2.795 0.350 3.125 1.010 ;
        RECT 3.355 0.085 3.685 0.820 ;
        RECT 4.355 0.085 4.615 1.010 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o41a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o41a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o41a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.528000 ;
    PORT
      LAYER li1 ;
        RECT 6.330 1.420 7.075 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.528000 ;
    PORT
      LAYER li1 ;
        RECT 7.805 0.505 8.035 0.670 ;
        RECT 7.305 0.335 8.035 0.505 ;
        RECT 7.305 0.255 7.635 0.335 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.528000 ;
    PORT
      LAYER li1 ;
        RECT 3.875 0.255 4.205 0.670 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.528000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.425 5.180 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 3.280 1.440 4.195 1.780 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.485 1.370 4.380 1.390 ;
        RECT 6.880 1.370 7.825 1.385 ;
        RECT 2.485 1.240 7.825 1.370 ;
        RECT 0.065 0.245 7.825 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.940 0.355 2.890 ;
        RECT 0.895 1.940 1.225 2.980 ;
        RECT 1.795 1.940 2.125 2.980 ;
        RECT 0.125 1.770 2.125 1.940 ;
        RECT 0.125 1.100 0.295 1.770 ;
        RECT 0.125 0.930 1.855 1.100 ;
        RECT 0.675 0.350 0.925 0.930 ;
        RECT 1.605 0.350 1.855 0.930 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.525 2.110 0.695 3.245 ;
        RECT 1.425 2.110 1.595 3.245 ;
        RECT 2.325 1.910 2.575 3.245 ;
        RECT 2.780 2.120 3.110 2.790 ;
        RECT 3.310 2.290 3.560 3.245 ;
        RECT 3.790 2.460 4.040 2.980 ;
        RECT 4.240 2.630 5.480 2.980 ;
        RECT 5.680 2.460 5.850 2.980 ;
        RECT 3.790 2.290 5.850 2.460 ;
        RECT 6.050 2.460 6.380 2.980 ;
        RECT 6.580 2.650 6.870 3.245 ;
        RECT 7.040 2.460 7.370 2.980 ;
        RECT 6.050 2.290 7.370 2.460 ;
        RECT 5.680 2.120 5.850 2.290 ;
        RECT 7.540 2.120 7.870 2.980 ;
        RECT 2.780 1.950 5.030 2.120 ;
        RECT 5.680 1.950 7.870 2.120 ;
        RECT 2.780 1.600 3.110 1.950 ;
        RECT 5.680 1.820 5.850 1.950 ;
        RECT 7.540 1.820 7.870 1.950 ;
        RECT 0.585 1.270 3.110 1.600 ;
        RECT 2.940 1.100 3.275 1.270 ;
        RECT 0.175 0.085 0.505 0.760 ;
        RECT 1.105 0.085 1.435 0.760 ;
        RECT 2.035 0.085 2.365 1.100 ;
        RECT 2.595 0.430 2.925 0.930 ;
        RECT 3.105 0.600 3.275 1.100 ;
        RECT 3.455 1.255 3.705 1.270 ;
        RECT 3.455 1.250 5.845 1.255 ;
        RECT 7.385 1.250 7.635 1.275 ;
        RECT 3.455 1.085 7.635 1.250 ;
        RECT 3.455 0.430 3.705 1.085 ;
        RECT 2.595 0.260 3.705 0.430 ;
        RECT 4.375 0.085 4.545 0.915 ;
        RECT 4.725 0.580 4.975 1.085 ;
        RECT 5.665 1.080 7.635 1.085 ;
        RECT 5.155 0.085 5.485 0.915 ;
        RECT 5.665 0.580 5.845 1.080 ;
        RECT 6.025 0.085 6.275 0.910 ;
        RECT 6.455 0.580 6.705 1.080 ;
        RECT 6.885 0.085 7.135 0.910 ;
        RECT 7.385 0.675 7.635 1.080 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__o41a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o41ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o41ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.810 1.350 3.235 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.920 2.295 2.890 ;
        RECT 2.125 1.680 2.295 1.920 ;
        RECT 2.125 1.350 2.525 1.680 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.680 1.795 2.890 ;
        RECT 1.565 1.350 1.955 1.680 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.350 1.385 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.220 0.245 3.330 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.602900 ;
    PORT
      LAYER li1 ;
        RECT 0.835 2.120 1.165 2.980 ;
        RECT 0.715 1.950 1.165 2.120 ;
        RECT 0.715 1.520 0.885 1.950 ;
        RECT 0.605 1.350 0.885 1.520 ;
        RECT 0.605 1.010 0.775 1.350 ;
        RECT 0.125 0.350 0.775 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.650 0.665 3.245 ;
        RECT 0.115 1.820 0.545 2.650 ;
        RECT 2.995 1.950 3.245 3.245 ;
        RECT 0.955 1.010 3.220 1.180 ;
        RECT 0.955 0.350 1.205 1.010 ;
        RECT 1.375 0.085 1.705 0.840 ;
        RECT 1.890 0.350 2.220 1.010 ;
        RECT 2.390 0.085 2.720 0.840 ;
        RECT 2.890 0.350 3.220 1.010 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o41ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o41ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o41ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 5.350 1.350 6.115 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.680 5.155 1.780 ;
        RECT 3.765 1.350 5.155 1.680 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 3.455 1.780 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.350 2.755 1.780 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.550 0.455 1.630 ;
        RECT 0.125 1.180 0.900 1.550 ;
        RECT 0.125 0.280 0.455 1.180 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.530 0.245 5.900 1.240 ;
        RECT 0.000 0.000 6.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.240 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.879200 ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.890 0.805 2.980 ;
        RECT 2.035 1.890 2.235 2.735 ;
        RECT 0.635 1.720 2.235 1.890 ;
        RECT 1.070 1.550 2.235 1.720 ;
        RECT 1.070 0.645 1.400 1.550 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.240 3.415 ;
        RECT 0.105 1.820 0.435 3.245 ;
        RECT 1.005 2.060 1.335 3.245 ;
        RECT 1.535 2.905 2.765 3.075 ;
        RECT 1.535 2.060 1.865 2.905 ;
        RECT 2.435 2.120 2.765 2.905 ;
        RECT 3.020 2.905 4.705 3.075 ;
        RECT 3.020 2.290 3.270 2.905 ;
        RECT 3.470 2.120 3.800 2.735 ;
        RECT 2.435 1.950 3.800 2.120 ;
        RECT 4.005 2.120 4.335 2.735 ;
        RECT 4.535 2.290 4.705 2.905 ;
        RECT 4.905 2.120 5.235 2.980 ;
        RECT 5.435 2.290 5.605 3.245 ;
        RECT 5.805 2.120 6.135 2.980 ;
        RECT 4.005 1.950 6.135 2.120 ;
        RECT 4.005 1.850 4.335 1.950 ;
        RECT 1.570 1.010 5.790 1.180 ;
        RECT 0.640 0.425 0.890 1.010 ;
        RECT 1.570 0.425 1.900 1.010 ;
        RECT 0.640 0.255 1.900 0.425 ;
        RECT 2.070 0.085 2.400 0.795 ;
        RECT 2.580 0.350 2.830 1.010 ;
        RECT 3.000 0.085 3.330 0.795 ;
        RECT 3.510 0.350 3.790 1.010 ;
        RECT 3.960 0.085 4.290 0.795 ;
        RECT 4.460 0.350 4.790 1.010 ;
        RECT 4.960 0.085 5.290 0.795 ;
        RECT 5.460 0.350 5.790 1.010 ;
        RECT 0.000 -0.085 6.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
  END
END sky130_fd_sc_hs__o41ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o41ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o41ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.180 9.955 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.180 8.035 1.550 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.395 1.180 6.115 1.550 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 3.160 1.550 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 1.145 1.550 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 10.075 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.586200 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.890 0.945 2.980 ;
        RECT 2.150 2.150 2.430 2.735 ;
        RECT 3.050 2.150 3.330 2.735 ;
        RECT 2.150 1.890 3.330 2.150 ;
        RECT 0.615 1.720 3.330 1.890 ;
        RECT 1.475 1.010 1.805 1.720 ;
        RECT 0.625 0.840 1.805 1.010 ;
        RECT 0.625 0.595 0.795 0.840 ;
        RECT 1.475 0.595 1.805 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.115 1.820 0.445 3.245 ;
        RECT 1.115 2.060 1.445 3.245 ;
        RECT 1.675 2.905 5.705 3.075 ;
        RECT 1.675 2.060 1.980 2.905 ;
        RECT 2.600 2.320 2.880 2.905 ;
        RECT 3.500 1.800 3.805 2.905 ;
        RECT 3.975 1.890 4.305 2.735 ;
        RECT 4.475 2.060 4.805 2.905 ;
        RECT 4.975 1.890 5.205 2.735 ;
        RECT 5.375 2.060 5.705 2.905 ;
        RECT 5.935 2.905 8.015 3.075 ;
        RECT 5.935 2.890 7.165 2.905 ;
        RECT 5.935 2.060 6.265 2.890 ;
        RECT 6.435 1.890 6.665 2.720 ;
        RECT 6.835 2.060 7.165 2.890 ;
        RECT 7.335 1.890 7.565 2.735 ;
        RECT 3.975 1.720 7.565 1.890 ;
        RECT 7.735 1.890 8.015 2.905 ;
        RECT 8.185 2.060 8.515 3.245 ;
        RECT 8.685 1.890 9.015 3.000 ;
        RECT 9.185 2.060 9.515 3.245 ;
        RECT 9.685 1.890 9.965 3.000 ;
        RECT 7.735 1.720 9.965 1.890 ;
        RECT 3.330 1.300 4.190 1.470 ;
        RECT 3.330 1.010 3.500 1.300 ;
        RECT 0.115 0.425 0.445 1.010 ;
        RECT 1.975 0.840 3.500 1.010 ;
        RECT 0.975 0.425 1.305 0.670 ;
        RECT 1.975 0.425 2.305 0.840 ;
        RECT 0.115 0.255 2.305 0.425 ;
        RECT 2.475 0.085 2.990 0.600 ;
        RECT 3.160 0.350 3.500 0.840 ;
        RECT 3.670 0.085 3.840 1.130 ;
        RECT 4.020 1.010 4.190 1.300 ;
        RECT 4.020 0.840 9.965 1.010 ;
        RECT 4.020 0.350 4.350 0.840 ;
        RECT 4.520 0.085 4.850 0.670 ;
        RECT 5.030 0.350 5.280 0.840 ;
        RECT 5.450 0.085 5.780 0.670 ;
        RECT 5.960 0.350 6.210 0.840 ;
        RECT 6.380 0.085 6.710 0.670 ;
        RECT 6.890 0.350 7.060 0.840 ;
        RECT 7.240 0.085 7.570 0.670 ;
        RECT 7.785 0.350 8.035 0.840 ;
        RECT 8.205 0.085 8.535 0.670 ;
        RECT 8.705 0.350 9.035 0.840 ;
        RECT 9.205 0.085 9.535 0.670 ;
        RECT 9.715 0.350 9.965 0.840 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__o41ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o211a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.335 1.470 2.005 1.800 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.255 3.715 0.640 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.490 3.335 1.800 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.635 1.490 4.195 1.800 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.155 1.240 4.245 1.450 ;
        RECT 0.005 0.245 4.245 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.820 0.445 2.980 ;
        RECT 0.085 1.130 0.255 1.820 ;
        RECT 0.085 0.350 0.445 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.615 2.310 1.855 3.245 ;
        RECT 2.395 2.140 2.725 2.980 ;
        RECT 2.895 2.310 3.705 3.245 ;
        RECT 3.875 2.140 4.205 2.980 ;
        RECT 0.925 1.970 4.205 2.140 ;
        RECT 0.925 1.650 1.095 1.970 ;
        RECT 2.395 1.940 2.835 1.970 ;
        RECT 0.425 1.320 1.095 1.650 ;
        RECT 2.665 1.320 2.835 1.940 ;
        RECT 1.265 1.130 2.495 1.300 ;
        RECT 2.665 1.150 4.135 1.320 ;
        RECT 0.615 0.085 0.945 1.130 ;
        RECT 1.265 0.660 1.595 1.130 ;
        RECT 2.325 0.980 2.495 1.130 ;
        RECT 1.765 0.085 2.155 0.925 ;
        RECT 2.325 0.810 3.185 0.980 ;
        RECT 3.760 0.835 4.135 1.150 ;
        RECT 3.885 0.660 4.135 0.835 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o211a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.350 2.295 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.335 1.350 1.795 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 1.125 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.820 3.225 2.980 ;
        RECT 3.005 1.410 3.225 1.820 ;
        RECT 3.005 1.130 3.235 1.410 ;
        RECT 2.980 0.350 3.235 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.105 2.120 0.435 2.860 ;
        RECT 0.605 2.290 0.935 3.245 ;
        RECT 1.105 2.120 1.435 2.860 ;
        RECT 2.025 2.290 2.725 3.245 ;
        RECT 0.105 1.950 2.675 2.120 ;
        RECT 0.105 1.820 0.435 1.950 ;
        RECT 2.505 1.630 2.675 1.950 ;
        RECT 3.395 1.820 3.725 3.245 ;
        RECT 2.505 1.300 2.835 1.630 ;
        RECT 2.505 1.180 2.675 1.300 ;
        RECT 0.605 1.010 2.675 1.180 ;
        RECT 0.130 0.350 0.775 1.010 ;
        RECT 1.025 0.670 2.350 0.840 ;
        RECT 1.025 0.350 1.355 0.670 ;
        RECT 1.525 0.085 1.775 0.500 ;
        RECT 2.020 0.350 2.350 0.670 ;
        RECT 2.550 0.085 2.800 0.840 ;
        RECT 3.410 0.085 3.740 1.130 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o211a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.075 1.450 6.595 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.450 5.835 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.435 2.835 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER li1 ;
        RECT 3.450 1.450 3.780 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.455 1.375 6.715 1.395 ;
        RECT 2.420 1.240 6.715 1.375 ;
        RECT 0.040 0.245 6.715 1.240 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.970 0.945 2.980 ;
        RECT 1.615 1.970 1.945 2.980 ;
        RECT 0.125 1.800 1.945 1.970 ;
        RECT 0.125 1.130 0.355 1.800 ;
        RECT 0.125 0.960 1.760 1.130 ;
        RECT 0.580 0.350 0.830 0.960 ;
        RECT 1.510 0.350 1.760 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.115 2.140 0.445 3.245 ;
        RECT 1.115 2.140 1.445 3.245 ;
        RECT 2.115 2.290 2.445 3.245 ;
        RECT 2.775 2.120 3.105 2.815 ;
        RECT 3.275 2.290 3.605 3.245 ;
        RECT 3.790 2.120 4.120 2.815 ;
        RECT 4.325 2.290 4.655 3.245 ;
        RECT 4.825 2.905 6.105 3.075 ;
        RECT 4.825 2.290 5.155 2.905 ;
        RECT 5.325 2.120 5.655 2.735 ;
        RECT 2.115 1.950 5.655 2.120 ;
        RECT 5.855 1.950 6.105 2.905 ;
        RECT 6.275 1.950 6.605 3.245 ;
        RECT 2.115 1.630 2.285 1.950 ;
        RECT 0.615 1.300 2.285 1.630 ;
        RECT 0.150 0.085 0.400 0.790 ;
        RECT 1.010 0.085 1.340 0.790 ;
        RECT 1.940 0.085 2.270 1.130 ;
        RECT 2.530 0.425 2.780 1.265 ;
        RECT 3.040 0.765 3.210 1.285 ;
        RECT 3.950 1.280 4.120 1.950 ;
        RECT 3.390 1.110 4.120 1.280 ;
        RECT 4.400 1.280 4.650 1.285 ;
        RECT 4.400 1.110 6.605 1.280 ;
        RECT 3.390 0.935 3.720 1.110 ;
        RECT 3.890 0.765 4.220 0.940 ;
        RECT 3.040 0.595 4.220 0.765 ;
        RECT 4.400 0.425 4.650 1.110 ;
        RECT 2.530 0.255 4.650 0.425 ;
        RECT 4.830 0.085 5.175 0.935 ;
        RECT 5.345 0.605 5.595 1.110 ;
        RECT 5.775 0.085 6.105 0.940 ;
        RECT 6.275 0.605 6.605 1.110 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__o211a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o211ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.630 0.835 2.890 ;
        RECT 0.605 1.550 1.165 1.630 ;
        RECT 0.665 1.300 1.165 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.405 1.300 1.795 1.630 ;
        RECT 1.565 0.440 1.795 1.300 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.180 2.305 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 2.875 1.240 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.427600 ;
    PORT
      LAYER li1 ;
        RECT 1.125 1.970 1.455 2.980 ;
        RECT 2.205 1.970 2.770 2.980 ;
        RECT 1.125 1.800 2.770 1.970 ;
        RECT 2.595 1.010 2.770 1.800 ;
        RECT 2.045 0.440 2.770 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.115 1.950 0.365 3.245 ;
        RECT 1.705 2.140 2.035 3.245 ;
        RECT 0.135 0.960 1.395 1.130 ;
        RECT 0.135 0.350 0.465 0.960 ;
        RECT 0.635 0.085 0.965 0.780 ;
        RECT 1.145 0.350 1.395 0.960 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__o211ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.685 1.320 4.695 1.650 ;
        RECT 4.365 1.180 4.695 1.320 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.650 3.235 1.780 ;
        RECT 2.435 1.320 3.445 1.650 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.350 2.015 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 1.240 2.440 1.290 ;
        RECT 0.020 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.215200 ;
    PORT
      LAYER li1 ;
        RECT 0.595 2.120 0.925 2.980 ;
        RECT 1.495 2.120 1.825 2.980 ;
        RECT 2.955 2.120 3.285 2.735 ;
        RECT 0.595 1.950 3.285 2.120 ;
        RECT 0.720 1.180 0.890 1.950 ;
        RECT 0.560 0.595 0.890 1.180 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.145 1.950 0.395 3.245 ;
        RECT 1.125 2.290 1.295 3.245 ;
        RECT 2.025 2.290 2.275 3.245 ;
        RECT 2.505 2.905 3.655 3.075 ;
        RECT 2.505 2.290 2.755 2.905 ;
        RECT 3.485 1.990 3.655 2.905 ;
        RECT 3.855 2.160 4.185 3.245 ;
        RECT 4.355 1.990 4.685 2.980 ;
        RECT 3.485 1.820 4.685 1.990 ;
        RECT 0.130 0.425 0.380 1.180 ;
        RECT 1.060 0.730 1.390 1.180 ;
        RECT 1.560 1.150 1.890 1.180 ;
        RECT 1.560 0.980 4.160 1.150 ;
        RECT 1.560 0.900 1.890 0.980 ;
        RECT 1.060 0.425 2.330 0.730 ;
        RECT 0.130 0.255 2.330 0.425 ;
        RECT 2.560 0.085 2.890 0.795 ;
        RECT 3.070 0.350 3.240 0.980 ;
        RECT 3.420 0.085 3.750 0.795 ;
        RECT 3.935 0.350 4.160 0.980 ;
        RECT 4.330 0.085 4.685 1.010 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o211ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.795 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 4.195 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 5.635 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 5.870 1.350 7.075 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.885 1.240 8.155 1.290 ;
        RECT 0.005 0.245 8.155 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.915200 ;
    PORT
      LAYER li1 ;
        RECT 2.430 2.120 2.760 2.735 ;
        RECT 3.380 2.120 3.710 2.735 ;
        RECT 4.940 2.120 5.270 2.980 ;
        RECT 5.940 2.120 6.270 2.980 ;
        RECT 7.545 2.120 8.035 2.890 ;
        RECT 2.430 1.950 8.035 2.120 ;
        RECT 7.365 1.550 8.035 1.950 ;
        RECT 7.365 1.180 7.545 1.550 ;
        RECT 6.505 1.010 7.545 1.180 ;
        RECT 6.505 0.595 6.675 1.010 ;
        RECT 7.365 0.595 7.545 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.130 2.120 0.460 2.980 ;
        RECT 0.660 2.290 0.830 3.245 ;
        RECT 1.030 2.120 1.360 2.980 ;
        RECT 1.560 2.290 1.730 3.245 ;
        RECT 1.930 2.905 4.210 3.075 ;
        RECT 1.930 2.120 2.260 2.905 ;
        RECT 2.960 2.290 3.210 2.905 ;
        RECT 3.880 2.290 4.210 2.905 ;
        RECT 4.440 2.290 4.770 3.245 ;
        RECT 5.440 2.290 5.770 3.245 ;
        RECT 6.440 2.290 7.290 3.245 ;
        RECT 0.130 1.950 2.260 2.120 ;
        RECT 0.115 1.010 5.765 1.180 ;
        RECT 0.115 0.350 0.445 1.010 ;
        RECT 0.615 0.085 0.945 0.840 ;
        RECT 1.125 0.350 1.375 1.010 ;
        RECT 1.545 0.085 1.875 0.840 ;
        RECT 2.055 0.350 2.225 1.010 ;
        RECT 2.405 0.085 2.735 0.840 ;
        RECT 2.915 0.350 3.085 1.010 ;
        RECT 3.265 0.085 3.595 0.840 ;
        RECT 3.795 0.820 4.905 1.010 ;
        RECT 3.795 0.350 3.965 0.820 ;
        RECT 5.085 0.650 5.255 0.840 ;
        RECT 4.145 0.425 5.255 0.650 ;
        RECT 5.435 0.595 5.765 1.010 ;
        RECT 5.995 0.425 6.325 1.180 ;
        RECT 6.855 0.425 7.185 0.840 ;
        RECT 7.715 0.425 8.045 1.180 ;
        RECT 4.145 0.255 8.045 0.425 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__o211ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o221a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.450 1.335 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.450 1.905 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.460 3.255 1.790 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.145 1.450 2.755 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.120 3.825 1.790 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 1.140 2.140 1.240 ;
        RECT 0.080 0.245 4.315 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.820 0.445 2.980 ;
        RECT 0.115 1.130 0.285 1.820 ;
        RECT 0.115 0.350 0.520 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.680 2.290 1.060 3.245 ;
        RECT 1.725 2.130 2.055 2.980 ;
        RECT 2.865 2.300 3.705 3.245 ;
        RECT 3.875 2.130 4.205 2.980 ;
        RECT 1.725 2.120 4.205 2.130 ;
        RECT 0.615 1.960 4.205 2.120 ;
        RECT 0.615 1.950 2.055 1.960 ;
        RECT 0.615 1.650 0.785 1.950 ;
        RECT 0.455 1.320 0.785 1.650 ;
        RECT 0.690 0.085 1.020 1.130 ;
        RECT 1.200 1.110 3.100 1.280 ;
        RECT 1.200 0.450 1.530 1.110 ;
        RECT 1.700 0.085 2.030 0.940 ;
        RECT 2.260 0.425 2.590 0.940 ;
        RECT 2.770 0.595 3.100 1.110 ;
        RECT 4.035 0.950 4.205 1.960 ;
        RECT 3.270 0.425 3.600 0.950 ;
        RECT 2.260 0.255 3.600 0.425 ;
        RECT 3.770 0.360 4.205 0.950 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o221a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.350 3.385 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.350 2.815 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.350 1.395 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.350 2.275 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.260 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.905 1.820 4.265 2.980 ;
        RECT 4.095 1.130 4.265 1.820 ;
        RECT 3.790 0.350 4.265 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 2.120 0.445 2.860 ;
        RECT 0.615 2.290 1.525 3.245 ;
        RECT 2.065 2.120 2.395 2.860 ;
        RECT 3.405 2.290 3.735 3.245 ;
        RECT 0.115 1.950 3.735 2.120 ;
        RECT 0.115 1.820 0.775 1.950 ;
        RECT 0.605 1.010 0.775 1.820 ;
        RECT 3.565 1.650 3.735 1.950 ;
        RECT 4.435 1.820 4.685 3.245 ;
        RECT 3.565 1.320 3.925 1.650 ;
        RECT 0.370 0.350 0.775 1.010 ;
        RECT 0.945 0.520 1.115 1.130 ;
        RECT 1.295 1.010 3.120 1.180 ;
        RECT 1.295 0.800 1.620 1.010 ;
        RECT 1.800 0.520 2.130 0.830 ;
        RECT 0.945 0.350 2.130 0.520 ;
        RECT 2.360 0.085 2.690 0.830 ;
        RECT 2.870 0.350 3.120 1.010 ;
        RECT 3.290 0.085 3.620 1.130 ;
        RECT 4.435 0.085 4.685 1.130 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o221a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.350 5.320 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.445 4.695 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.445 4.195 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.445 2.755 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.445 0.890 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.365 3.280 1.395 ;
        RECT 0.005 0.245 7.675 1.365 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.235700 ;
    PORT
      LAYER li1 ;
        RECT 5.830 2.020 6.160 2.980 ;
        RECT 6.785 2.020 7.115 2.980 ;
        RECT 5.830 1.850 7.115 2.020 ;
        RECT 6.785 1.780 7.115 1.850 ;
        RECT 6.785 1.550 7.555 1.780 ;
        RECT 6.785 1.180 7.065 1.550 ;
        RECT 5.735 1.010 7.065 1.180 ;
        RECT 5.735 0.475 5.985 1.010 ;
        RECT 6.735 0.475 7.065 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.115 1.950 0.365 3.245 ;
        RECT 0.565 2.120 0.895 2.955 ;
        RECT 1.095 2.290 1.345 3.245 ;
        RECT 1.515 2.905 2.745 3.075 ;
        RECT 1.515 2.290 1.845 2.905 ;
        RECT 2.045 2.120 2.215 2.735 ;
        RECT 2.415 2.290 2.745 2.905 ;
        RECT 2.915 2.290 3.630 3.245 ;
        RECT 3.800 2.905 5.130 3.075 ;
        RECT 3.800 2.290 4.130 2.905 ;
        RECT 4.300 2.120 4.630 2.735 ;
        RECT 4.800 2.290 5.130 2.905 ;
        RECT 5.300 2.290 5.630 3.245 ;
        RECT 6.360 2.190 6.610 3.245 ;
        RECT 0.565 1.950 5.660 2.120 ;
        RECT 7.315 1.950 7.565 3.245 ;
        RECT 1.060 1.275 1.230 1.950 ;
        RECT 5.490 1.680 5.660 1.950 ;
        RECT 5.490 1.350 6.615 1.680 ;
        RECT 0.115 0.435 0.365 1.275 ;
        RECT 0.545 1.105 1.230 1.275 ;
        RECT 1.475 1.275 1.805 1.285 ;
        RECT 1.475 1.180 4.115 1.275 ;
        RECT 1.475 1.105 5.055 1.180 ;
        RECT 0.545 0.605 0.795 1.105 ;
        RECT 1.475 1.025 2.740 1.105 ;
        RECT 0.975 0.435 1.305 0.935 ;
        RECT 1.475 0.605 1.805 1.025 ;
        RECT 1.975 0.455 2.305 0.855 ;
        RECT 2.475 0.635 2.670 1.025 ;
        RECT 3.940 1.010 5.055 1.105 ;
        RECT 2.840 0.455 3.170 0.855 ;
        RECT 1.975 0.435 3.170 0.455 ;
        RECT 0.115 0.285 3.170 0.435 ;
        RECT 0.115 0.265 2.305 0.285 ;
        RECT 3.430 0.085 3.760 0.935 ;
        RECT 3.940 0.585 4.115 1.010 ;
        RECT 4.295 0.085 4.625 0.840 ;
        RECT 4.805 0.590 5.055 1.010 ;
        RECT 5.235 0.085 5.565 1.180 ;
        RECT 6.165 0.085 6.565 0.805 ;
        RECT 7.235 0.085 7.565 1.255 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__o221a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.300 3.715 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.680 2.775 2.890 ;
        RECT 2.445 1.350 2.775 1.680 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.350 1.635 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.875 1.350 2.275 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.835 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.011700 ;
    PORT
      LAYER li1 ;
        RECT 0.325 2.120 0.575 2.980 ;
        RECT 2.025 2.120 2.355 2.980 ;
        RECT 0.325 1.950 2.355 2.120 ;
        RECT 0.605 1.130 0.775 1.950 ;
        RECT 0.115 0.960 0.775 1.130 ;
        RECT 0.115 0.350 0.445 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.745 2.290 1.560 3.245 ;
        RECT 3.165 1.950 3.495 3.245 ;
        RECT 1.175 1.130 2.505 1.180 ;
        RECT 1.175 1.010 3.725 1.130 ;
        RECT 1.175 0.800 1.505 1.010 ;
        RECT 2.175 0.960 3.725 1.010 ;
        RECT 0.615 0.520 0.945 0.770 ;
        RECT 1.675 0.520 2.005 0.795 ;
        RECT 0.615 0.350 2.005 0.520 ;
        RECT 2.175 0.350 2.505 0.960 ;
        RECT 2.675 0.085 3.225 0.790 ;
        RECT 3.395 0.350 3.725 0.960 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o221ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.645 1.950 5.635 2.120 ;
        RECT 3.645 1.350 3.975 1.950 ;
        RECT 4.925 1.350 5.635 1.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.345 1.350 4.675 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.950 3.405 2.120 ;
        RECT 1.085 1.350 2.275 1.950 ;
        RECT 3.075 1.350 3.405 1.950 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.520 1.350 2.850 1.780 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.425 1.240 5.755 1.295 ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.232000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 2.460 0.855 2.980 ;
        RECT 2.365 2.460 2.695 2.735 ;
        RECT 4.365 2.460 4.615 2.735 ;
        RECT 0.605 2.290 4.615 2.460 ;
        RECT 0.605 0.595 0.875 2.290 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.155 1.950 0.405 3.245 ;
        RECT 1.055 2.630 1.695 3.245 ;
        RECT 1.865 2.905 3.195 3.075 ;
        RECT 1.865 2.630 2.195 2.905 ;
        RECT 2.865 2.630 3.195 2.905 ;
        RECT 3.365 2.630 3.695 3.245 ;
        RECT 3.865 2.905 5.145 3.075 ;
        RECT 3.865 2.630 4.195 2.905 ;
        RECT 4.815 2.290 5.145 2.905 ;
        RECT 5.315 2.290 5.645 3.245 ;
        RECT 0.115 0.425 0.365 1.130 ;
        RECT 1.055 1.010 3.280 1.180 ;
        RECT 1.055 0.425 1.305 1.010 ;
        RECT 0.115 0.255 1.305 0.425 ;
        RECT 1.535 0.425 1.865 0.820 ;
        RECT 2.045 0.595 2.215 1.010 ;
        RECT 2.395 0.425 2.725 0.820 ;
        RECT 2.895 0.595 3.280 1.010 ;
        RECT 3.460 1.010 5.645 1.180 ;
        RECT 3.460 0.425 3.710 1.010 ;
        RECT 1.535 0.255 3.710 0.425 ;
        RECT 3.880 0.085 4.210 0.820 ;
        RECT 4.380 0.405 4.710 1.010 ;
        RECT 4.880 0.085 5.210 0.820 ;
        RECT 5.390 0.405 5.645 1.010 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__o221ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o221ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.210 1.260 6.575 1.590 ;
        RECT 8.285 1.260 9.955 1.780 ;
        RECT 6.405 1.090 8.455 1.260 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.430 8.035 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.710 6.000 1.880 ;
        RECT 2.545 1.350 3.555 1.710 ;
        RECT 5.405 1.350 6.000 1.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 4.185 1.180 5.195 1.540 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.405 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 2.275 1.290 ;
        RECT 0.005 0.245 10.075 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.514400 ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.120 0.895 2.980 ;
        RECT 1.575 2.220 1.825 2.980 ;
        RECT 4.055 2.220 4.225 2.735 ;
        RECT 4.925 2.220 5.255 2.735 ;
        RECT 6.930 2.520 7.260 2.735 ;
        RECT 6.845 2.220 7.260 2.520 ;
        RECT 1.575 2.120 7.260 2.220 ;
        RECT 7.830 2.120 8.160 2.735 ;
        RECT 0.565 2.050 8.160 2.120 ;
        RECT 0.565 1.950 1.825 2.050 ;
        RECT 6.845 1.950 8.160 2.050 ;
        RECT 1.575 1.820 1.825 1.950 ;
        RECT 1.575 1.180 1.745 1.820 ;
        RECT 0.545 1.010 1.745 1.180 ;
        RECT 0.545 0.595 0.875 1.010 ;
        RECT 1.405 0.595 1.745 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.115 1.950 0.365 3.245 ;
        RECT 1.065 2.290 1.395 3.245 ;
        RECT 2.025 2.390 2.355 3.245 ;
        RECT 2.525 2.560 2.855 2.980 ;
        RECT 3.025 2.730 3.355 3.245 ;
        RECT 3.525 2.905 5.755 3.075 ;
        RECT 3.525 2.560 3.855 2.905 ;
        RECT 2.525 2.390 3.855 2.560 ;
        RECT 4.425 2.390 4.755 2.905 ;
        RECT 5.425 2.390 5.755 2.905 ;
        RECT 5.925 2.390 6.255 3.245 ;
        RECT 6.425 2.905 8.530 3.075 ;
        RECT 6.425 2.730 6.760 2.905 ;
        RECT 6.425 2.650 6.675 2.730 ;
        RECT 7.460 2.290 7.630 2.905 ;
        RECT 8.360 2.120 8.530 2.905 ;
        RECT 8.730 2.290 8.980 3.245 ;
        RECT 9.180 2.120 9.510 2.980 ;
        RECT 8.360 1.950 9.510 2.120 ;
        RECT 9.710 1.950 9.960 3.245 ;
        RECT 0.115 0.425 0.375 1.180 ;
        RECT 1.915 1.010 4.015 1.180 ;
        RECT 5.405 1.010 5.735 1.050 ;
        RECT 1.045 0.425 1.235 0.840 ;
        RECT 1.915 0.770 3.155 1.010 ;
        RECT 1.915 0.425 2.165 0.770 ;
        RECT 3.335 0.600 3.505 0.840 ;
        RECT 3.685 0.770 5.735 1.010 ;
        RECT 5.905 0.920 6.235 1.090 ;
        RECT 8.775 0.920 9.965 1.090 ;
        RECT 5.905 0.750 9.025 0.920 ;
        RECT 5.905 0.600 6.235 0.750 ;
        RECT 0.115 0.255 2.165 0.425 ;
        RECT 2.395 0.350 6.235 0.600 ;
        RECT 6.405 0.085 6.735 0.580 ;
        RECT 6.905 0.350 7.155 0.750 ;
        RECT 7.335 0.085 7.665 0.580 ;
        RECT 7.835 0.350 8.085 0.750 ;
        RECT 8.265 0.085 8.605 0.580 ;
        RECT 8.775 0.350 9.025 0.750 ;
        RECT 9.205 0.085 9.535 0.750 ;
        RECT 9.715 0.350 9.965 0.920 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__o221ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o311a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o311a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.015 1.120 3.385 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.635 2.320 2.845 2.490 ;
        RECT 1.635 1.470 1.805 2.320 ;
        RECT 1.455 1.140 1.805 1.470 ;
        RECT 2.515 1.445 2.845 2.320 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.120 2.305 2.150 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.920 1.140 1.285 1.470 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.140 0.410 1.470 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.365 1.140 4.310 1.240 ;
        RECT 0.090 0.245 4.310 1.140 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.960 4.235 2.980 ;
        RECT 4.065 1.130 4.235 1.960 ;
        RECT 3.870 0.350 4.235 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.135 1.810 0.465 2.955 ;
        RECT 0.635 1.980 0.965 3.245 ;
        RECT 1.135 2.785 3.185 2.955 ;
        RECT 1.135 1.810 1.465 2.785 ;
        RECT 0.135 1.640 1.465 1.810 ;
        RECT 3.015 1.790 3.185 2.785 ;
        RECT 3.355 1.960 3.685 3.245 ;
        RECT 0.580 0.970 0.750 1.640 ;
        RECT 3.015 1.620 3.895 1.790 ;
        RECT 3.595 1.350 3.895 1.620 ;
        RECT 0.200 0.800 0.750 0.970 ;
        RECT 0.200 0.350 0.530 0.800 ;
        RECT 1.060 0.610 1.390 0.970 ;
        RECT 1.560 0.780 3.690 0.950 ;
        RECT 1.060 0.280 3.180 0.610 ;
        RECT 3.360 0.085 3.690 0.780 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o311a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o311a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o311a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 2.925 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.350 2.355 2.890 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.350 1.815 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.350 1.315 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.330 1.890 3.660 2.980 ;
        RECT 3.330 1.720 4.195 1.890 ;
        RECT 3.965 1.050 4.195 1.720 ;
        RECT 3.435 0.810 4.195 1.050 ;
        RECT 3.435 0.350 3.685 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.225 2.120 0.605 2.860 ;
        RECT 0.775 2.290 1.105 3.245 ;
        RECT 1.335 2.120 1.665 2.980 ;
        RECT 0.225 1.950 1.665 2.120 ;
        RECT 2.745 1.950 3.075 3.245 ;
        RECT 3.830 2.060 4.160 3.245 ;
        RECT 0.225 1.820 0.775 1.950 ;
        RECT 0.605 1.180 0.775 1.820 ;
        RECT 3.095 1.220 3.510 1.550 ;
        RECT 3.095 1.180 3.265 1.220 ;
        RECT 0.605 1.010 3.265 1.180 ;
        RECT 0.205 0.350 0.775 1.010 ;
        RECT 1.180 0.670 2.660 0.840 ;
        RECT 1.180 0.350 1.510 0.670 ;
        RECT 1.690 0.085 2.150 0.500 ;
        RECT 2.330 0.350 2.660 0.670 ;
        RECT 2.830 0.085 3.160 0.840 ;
        RECT 3.855 0.085 4.205 0.600 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__o311a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o311a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o311a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 7.105 1.470 8.035 1.800 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 6.525 1.300 6.935 1.550 ;
        RECT 8.205 1.300 8.535 1.780 ;
        RECT 6.525 1.220 8.535 1.300 ;
        RECT 6.765 1.130 8.535 1.220 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.870 1.420 6.200 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.640 5.360 1.800 ;
        RECT 2.505 1.265 2.910 1.550 ;
        RECT 3.995 1.470 5.360 1.640 ;
        RECT 3.995 1.265 4.165 1.470 ;
        RECT 2.505 1.220 4.165 1.265 ;
        RECT 2.740 1.095 4.165 1.220 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.435 3.825 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.160 2.680 1.240 ;
        RECT 4.145 1.160 4.695 1.375 ;
        RECT 0.005 0.245 8.635 1.160 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.345400 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.890 0.895 2.980 ;
        RECT 1.565 1.890 1.895 2.980 ;
        RECT 0.565 1.720 1.895 1.890 ;
        RECT 0.565 1.650 0.895 1.720 ;
        RECT 0.125 1.480 0.895 1.650 ;
        RECT 0.125 1.310 0.355 1.480 ;
        RECT 0.125 1.140 0.945 1.310 ;
        RECT 0.615 1.050 0.945 1.140 ;
        RECT 0.615 0.880 2.070 1.050 ;
        RECT 0.615 0.350 0.945 0.880 ;
        RECT 1.740 0.350 2.070 0.880 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 1.065 2.060 1.395 3.245 ;
        RECT 2.150 2.060 2.480 3.245 ;
        RECT 2.655 2.120 2.985 2.980 ;
        RECT 3.225 2.290 3.920 3.245 ;
        RECT 4.090 2.140 4.420 2.980 ;
        RECT 4.590 2.540 4.920 3.245 ;
        RECT 6.220 2.960 8.525 3.075 ;
        RECT 5.150 2.905 8.525 2.960 ;
        RECT 5.150 2.710 6.550 2.905 ;
        RECT 6.720 2.565 8.025 2.735 ;
        RECT 4.590 2.395 6.550 2.540 ;
        RECT 4.590 2.370 7.575 2.395 ;
        RECT 4.590 2.310 4.920 2.370 ;
        RECT 5.750 2.140 6.100 2.200 ;
        RECT 4.090 2.120 6.100 2.140 ;
        RECT 2.655 1.970 6.100 2.120 ;
        RECT 6.380 1.970 7.575 2.370 ;
        RECT 7.775 1.970 8.025 2.565 ;
        RECT 8.195 1.970 8.525 2.905 ;
        RECT 2.655 1.950 4.420 1.970 ;
        RECT 2.655 1.890 2.985 1.950 ;
        RECT 4.090 1.940 4.420 1.950 ;
        RECT 5.530 1.950 6.100 1.970 ;
        RECT 2.095 1.720 2.985 1.890 ;
        RECT 2.095 1.550 2.265 1.720 ;
        RECT 1.255 1.220 2.265 1.550 ;
        RECT 5.530 1.300 5.700 1.950 ;
        RECT 4.335 1.130 5.700 1.300 ;
        RECT 0.115 0.085 0.445 0.970 ;
        RECT 1.115 0.085 1.570 0.680 ;
        RECT 2.240 0.085 2.570 1.050 ;
        RECT 4.335 0.935 4.585 1.130 ;
        RECT 6.265 0.960 6.595 1.050 ;
        RECT 2.800 0.425 3.130 0.925 ;
        RECT 3.300 0.765 4.075 0.925 ;
        RECT 4.765 0.765 5.095 0.960 ;
        RECT 3.300 0.595 5.095 0.765 ;
        RECT 5.265 0.790 8.525 0.960 ;
        RECT 5.265 0.425 5.595 0.790 ;
        RECT 2.800 0.255 5.595 0.425 ;
        RECT 5.765 0.085 6.095 0.620 ;
        RECT 6.265 0.370 6.595 0.790 ;
        RECT 6.765 0.085 7.095 0.620 ;
        RECT 7.265 0.350 7.595 0.790 ;
        RECT 7.765 0.085 8.095 0.620 ;
        RECT 8.275 0.350 8.525 0.790 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__o311a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o311ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o311ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.705 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.350 1.315 2.890 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.180 1.845 1.550 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.180 2.415 1.550 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.180 3.255 1.550 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.220 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.011700 ;
    PORT
      LAYER li1 ;
        RECT 1.785 1.890 2.115 2.980 ;
        RECT 2.805 1.890 3.235 2.980 ;
        RECT 1.785 1.720 3.235 1.890 ;
        RECT 2.585 1.010 2.755 1.720 ;
        RECT 2.585 0.350 3.110 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.225 1.950 0.555 3.245 ;
        RECT 2.285 2.060 2.615 3.245 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 0.615 1.010 0.945 1.130 ;
        RECT 0.615 0.840 2.220 1.010 ;
        RECT 0.615 0.350 0.945 0.840 ;
        RECT 1.115 0.085 1.675 0.650 ;
        RECT 1.890 0.330 2.220 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o311ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o311ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o311ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.835 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.350 2.275 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 3.235 1.780 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 4.195 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.300 5.635 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.754600 ;
    PORT
      LAYER li1 ;
        RECT 2.600 2.120 2.930 2.735 ;
        RECT 3.500 2.120 3.750 2.980 ;
        RECT 4.480 2.120 4.650 2.980 ;
        RECT 5.300 2.120 5.630 2.980 ;
        RECT 2.600 1.950 5.630 2.120 ;
        RECT 4.400 1.130 4.730 1.950 ;
        RECT 4.400 0.960 5.645 1.130 ;
        RECT 4.400 0.595 4.705 0.960 ;
        RECT 5.395 0.350 5.645 0.960 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.120 2.120 0.450 2.980 ;
        RECT 0.650 2.290 0.900 3.245 ;
        RECT 1.070 2.120 1.400 2.980 ;
        RECT 1.590 2.905 3.300 3.075 ;
        RECT 1.590 2.290 1.920 2.905 ;
        RECT 2.120 2.120 2.370 2.735 ;
        RECT 3.130 2.290 3.300 2.905 ;
        RECT 3.950 2.290 4.280 3.245 ;
        RECT 4.850 2.290 5.100 3.245 ;
        RECT 0.120 1.950 2.370 2.120 ;
        RECT 0.115 1.010 4.225 1.180 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.840 ;
        RECT 1.115 0.350 1.365 1.010 ;
        RECT 1.535 0.085 1.865 0.840 ;
        RECT 2.045 0.350 2.295 1.010 ;
        RECT 2.465 0.085 2.795 0.840 ;
        RECT 2.975 0.350 3.225 1.010 ;
        RECT 3.395 0.425 3.725 0.840 ;
        RECT 3.895 0.595 4.225 1.010 ;
        RECT 4.885 0.425 5.215 0.790 ;
        RECT 3.395 0.255 5.215 0.425 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__o311ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o311ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o311ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 9.165 1.350 10.435 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.350 7.775 1.780 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 5.185 1.640 6.195 1.780 ;
        RECT 4.485 1.430 6.195 1.640 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 2.245 1.430 4.195 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 1.240 1.780 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 11.035 1.240 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.271700 ;
    PORT
      LAYER li1 ;
        RECT 0.740 2.120 1.070 2.980 ;
        RECT 1.740 2.120 2.070 2.980 ;
        RECT 4.685 2.120 5.015 2.735 ;
        RECT 5.685 2.120 6.015 2.735 ;
        RECT 0.740 1.950 6.595 2.120 ;
        RECT 1.740 1.820 2.070 1.950 ;
        RECT 4.685 1.820 5.015 1.950 ;
        RECT 6.365 1.260 6.595 1.950 ;
        RECT 1.410 1.100 6.595 1.260 ;
        RECT 0.545 1.090 6.595 1.100 ;
        RECT 0.545 0.770 1.740 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.115 1.950 0.445 3.245 ;
        RECT 1.240 2.290 1.570 3.245 ;
        RECT 2.240 2.290 3.905 3.245 ;
        RECT 4.185 2.905 8.565 3.075 ;
        RECT 4.185 2.290 4.515 2.905 ;
        RECT 5.185 2.290 5.515 2.905 ;
        RECT 6.285 2.290 6.615 2.905 ;
        RECT 6.785 2.120 7.115 2.735 ;
        RECT 7.285 2.290 7.615 2.905 ;
        RECT 7.785 2.150 8.065 2.735 ;
        RECT 8.235 2.330 8.565 2.905 ;
        RECT 8.795 2.330 9.125 3.245 ;
        RECT 9.295 2.150 9.525 2.980 ;
        RECT 9.695 2.330 10.025 3.245 ;
        RECT 10.195 2.150 10.475 2.980 ;
        RECT 7.785 2.120 10.475 2.150 ;
        RECT 6.785 1.950 10.475 2.120 ;
        RECT 10.675 1.820 10.925 3.245 ;
        RECT 7.945 1.300 8.975 1.470 ;
        RECT 7.945 1.180 8.115 1.300 ;
        RECT 0.115 0.600 0.365 1.130 ;
        RECT 6.890 1.010 8.115 1.180 ;
        RECT 8.725 1.130 8.975 1.300 ;
        RECT 6.890 0.920 7.140 1.010 ;
        RECT 1.920 0.750 3.900 0.920 ;
        RECT 4.070 0.750 7.140 0.920 ;
        RECT 1.920 0.600 2.090 0.750 ;
        RECT 0.115 0.350 2.090 0.600 ;
        RECT 4.070 0.580 4.240 0.750 ;
        RECT 2.270 0.330 4.240 0.580 ;
        RECT 4.410 0.085 4.740 0.580 ;
        RECT 4.920 0.350 5.170 0.750 ;
        RECT 5.350 0.085 5.680 0.580 ;
        RECT 5.860 0.350 6.190 0.750 ;
        RECT 6.370 0.085 6.710 0.580 ;
        RECT 6.890 0.350 7.140 0.750 ;
        RECT 7.320 0.085 7.650 0.825 ;
        RECT 7.945 0.350 8.115 1.010 ;
        RECT 8.295 0.085 8.545 1.130 ;
        RECT 8.725 0.960 10.415 1.130 ;
        RECT 8.725 0.350 8.975 0.960 ;
        RECT 9.155 0.085 9.995 0.790 ;
        RECT 10.165 0.350 10.415 0.960 ;
        RECT 10.595 0.085 10.925 1.130 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__o311ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o2111a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2111a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.300 3.735 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.715 1.415 3.235 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.415 2.505 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 0.440 1.875 1.900 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.550 1.335 1.880 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.820 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.533900 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.820 0.445 2.980 ;
        RECT 0.095 1.040 0.265 1.820 ;
        RECT 0.095 0.350 0.355 1.040 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.615 2.410 0.945 3.245 ;
        RECT 1.195 2.245 1.525 2.925 ;
        RECT 1.740 2.455 2.290 3.245 ;
        RECT 2.535 2.245 2.865 2.925 ;
        RECT 1.195 2.240 2.865 2.245 ;
        RECT 0.615 2.070 2.865 2.240 ;
        RECT 0.615 1.550 0.785 2.070 ;
        RECT 2.535 2.045 2.865 2.070 ;
        RECT 3.405 1.950 3.735 3.245 ;
        RECT 0.435 1.380 0.785 1.550 ;
        RECT 0.435 1.210 1.330 1.380 ;
        RECT 0.535 0.085 0.865 1.040 ;
        RECT 1.080 0.350 1.330 1.210 ;
        RECT 2.380 0.960 3.710 1.130 ;
        RECT 2.380 0.350 2.710 0.960 ;
        RECT 2.880 0.085 3.210 0.790 ;
        RECT 3.380 0.350 3.710 0.960 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__o2111a_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o2111a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2111a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.835 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.180 1.345 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.180 1.915 1.550 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.155 1.350 2.755 1.780 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.261000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.350 3.255 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 0.245 4.795 1.240 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.820 4.185 2.980 ;
        RECT 4.015 1.130 4.185 1.820 ;
        RECT 3.910 0.350 4.240 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.295 1.820 0.625 3.245 ;
        RECT 1.285 2.120 1.615 2.860 ;
        RECT 1.785 2.290 2.115 3.245 ;
        RECT 2.375 2.120 2.705 2.880 ;
        RECT 2.875 2.290 3.685 3.245 ;
        RECT 1.285 1.950 3.685 2.120 ;
        RECT 1.285 1.820 1.615 1.950 ;
        RECT 3.515 1.630 3.685 1.950 ;
        RECT 4.355 1.820 4.685 3.245 ;
        RECT 3.515 1.300 3.845 1.630 ;
        RECT 3.515 1.180 3.685 1.300 ;
        RECT 2.850 1.010 3.685 1.180 ;
        RECT 0.250 0.840 1.720 1.010 ;
        RECT 0.250 0.350 0.580 0.840 ;
        RECT 0.750 0.085 1.220 0.670 ;
        RECT 1.390 0.350 1.720 0.840 ;
        RECT 2.850 0.350 3.180 1.010 ;
        RECT 3.410 0.085 3.740 0.825 ;
        RECT 4.420 0.085 4.685 1.130 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__o2111a_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o2111a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2111a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 5.325 1.450 5.655 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.522000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.450 5.155 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.474000 ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.450 3.315 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.474000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.450 1.795 1.780 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.474000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.550 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.255 1.240 4.675 1.410 ;
        RECT 0.005 0.245 8.125 1.240 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.142400 ;
    PORT
      LAYER li1 ;
        RECT 6.315 2.180 6.590 2.980 ;
        RECT 7.295 2.180 7.545 2.980 ;
        RECT 6.315 1.850 7.545 2.180 ;
        RECT 7.295 1.650 7.545 1.850 ;
        RECT 7.295 1.480 8.035 1.650 ;
        RECT 7.805 1.180 8.035 1.480 ;
        RECT 6.185 1.010 8.035 1.180 ;
        RECT 6.185 0.350 6.515 1.010 ;
        RECT 7.185 0.350 7.515 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.115 2.120 0.445 2.820 ;
        RECT 0.615 2.315 0.945 3.245 ;
        RECT 1.115 2.120 1.445 2.820 ;
        RECT 1.615 2.315 1.945 3.245 ;
        RECT 2.150 2.120 2.480 2.820 ;
        RECT 2.685 2.315 3.015 3.245 ;
        RECT 3.220 2.905 4.550 3.075 ;
        RECT 3.220 2.120 3.550 2.905 ;
        RECT 3.720 2.460 4.050 2.735 ;
        RECT 4.220 2.630 4.550 2.905 ;
        RECT 4.780 2.630 5.110 3.245 ;
        RECT 5.280 2.460 5.610 2.980 ;
        RECT 3.720 2.290 5.610 2.460 ;
        RECT 5.815 2.290 6.145 3.245 ;
        RECT 6.765 2.350 7.095 3.245 ;
        RECT 0.115 1.950 6.145 2.120 ;
        RECT 0.720 1.130 0.890 1.950 ;
        RECT 2.150 1.940 2.480 1.950 ;
        RECT 5.975 1.680 6.145 1.950 ;
        RECT 7.715 1.820 8.045 3.245 ;
        RECT 5.975 1.350 7.125 1.680 ;
        RECT 2.365 1.280 2.775 1.300 ;
        RECT 0.115 0.600 0.380 1.115 ;
        RECT 0.550 0.770 0.890 1.130 ;
        RECT 1.060 0.600 1.230 1.130 ;
        RECT 0.115 0.425 1.230 0.600 ;
        RECT 1.410 0.880 1.740 1.130 ;
        RECT 2.365 1.110 5.505 1.280 ;
        RECT 2.365 1.050 3.555 1.110 ;
        RECT 1.410 0.710 3.125 0.880 ;
        RECT 1.410 0.595 1.740 0.710 ;
        RECT 1.920 0.425 2.250 0.540 ;
        RECT 2.875 0.520 3.125 0.710 ;
        RECT 3.305 0.520 3.555 1.050 ;
        RECT 0.115 0.255 2.250 0.425 ;
        RECT 3.735 0.085 4.065 0.940 ;
        RECT 4.235 0.520 4.565 1.110 ;
        RECT 4.825 0.085 5.155 0.940 ;
        RECT 5.335 0.350 5.505 1.110 ;
        RECT 5.685 0.085 6.015 1.130 ;
        RECT 6.685 0.085 7.015 0.815 ;
        RECT 7.685 0.085 8.015 0.815 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__o2111a_4

#--------EOF---------

MACRO sky130_fd_sc_hs__o2111ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2111ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.180 3.255 1.550 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 2.200 1.180 2.755 1.550 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.595 1.180 1.990 1.550 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.440 1.425 1.550 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.180 0.910 1.550 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.355 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.162500 ;
    PORT
      LAYER li1 ;
        RECT 0.880 1.890 1.315 2.980 ;
        RECT 1.985 1.890 2.315 2.980 ;
        RECT 0.115 1.720 2.315 1.890 ;
        RECT 0.115 1.010 0.285 1.720 ;
        RECT 0.115 0.350 0.785 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.380 2.060 0.710 3.245 ;
        RECT 1.485 2.060 1.815 3.245 ;
        RECT 2.890 1.820 3.220 3.245 ;
        RECT 1.825 0.840 3.245 1.010 ;
        RECT 1.825 0.350 2.155 0.840 ;
        RECT 2.325 0.085 2.745 0.600 ;
        RECT 2.915 0.350 3.245 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__o2111ai_1

#--------EOF---------

MACRO sky130_fd_sc_hs__o2111ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2111ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.350 5.635 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.350 4.675 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.350 3.715 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 1.345 1.300 2.015 1.630 ;
        RECT 1.565 1.180 1.795 1.300 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.245 5.710 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.551200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.970 0.935 2.980 ;
        RECT 1.555 2.120 1.885 2.980 ;
        RECT 2.455 2.120 2.785 2.980 ;
        RECT 3.915 2.120 4.245 2.735 ;
        RECT 1.555 1.970 4.245 2.120 ;
        RECT 0.605 1.950 4.245 1.970 ;
        RECT 0.605 1.800 1.885 1.950 ;
        RECT 0.605 1.180 0.935 1.800 ;
        RECT 0.690 1.130 0.935 1.180 ;
        RECT 0.690 0.595 0.940 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.155 1.820 0.405 3.245 ;
        RECT 1.105 2.140 1.355 3.245 ;
        RECT 2.085 2.290 2.255 3.245 ;
        RECT 2.985 2.290 3.235 3.245 ;
        RECT 3.465 2.905 4.615 3.075 ;
        RECT 3.465 2.290 3.715 2.905 ;
        RECT 4.445 2.120 4.615 2.905 ;
        RECT 4.815 2.290 5.145 3.245 ;
        RECT 5.315 2.120 5.645 2.980 ;
        RECT 4.445 1.950 5.645 2.120 ;
        RECT 1.120 1.010 1.290 1.130 ;
        RECT 1.970 1.010 2.300 1.130 ;
        RECT 0.180 0.425 0.510 1.010 ;
        RECT 1.120 0.840 2.300 1.010 ;
        RECT 1.120 0.425 1.290 0.840 ;
        RECT 0.180 0.255 1.290 0.425 ;
        RECT 1.470 0.425 1.800 0.670 ;
        RECT 1.970 0.595 2.300 0.840 ;
        RECT 2.530 1.010 5.600 1.180 ;
        RECT 2.530 0.595 2.860 1.010 ;
        RECT 3.030 0.425 3.360 0.840 ;
        RECT 1.470 0.255 3.360 0.425 ;
        RECT 3.540 0.350 3.710 1.010 ;
        RECT 3.890 0.085 4.220 0.840 ;
        RECT 4.420 0.350 4.670 1.010 ;
        RECT 4.840 0.085 5.170 0.840 ;
        RECT 5.350 0.350 5.600 1.010 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__o2111ai_2

#--------EOF---------

MACRO sky130_fd_sc_hs__o2111ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o2111ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 6.285 1.350 7.635 1.780 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.350 9.490 1.780 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.350 6.115 1.780 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.630 4.195 1.780 ;
        RECT 2.210 1.300 4.195 1.630 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 1.350 1.780 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 10.075 1.240 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.411800 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.120 1.200 2.980 ;
        RECT 1.870 2.120 2.200 2.980 ;
        RECT 0.115 1.970 2.200 2.120 ;
        RECT 3.190 2.120 3.520 2.980 ;
        RECT 4.190 2.120 4.520 2.980 ;
        RECT 8.185 2.120 8.515 2.735 ;
        RECT 9.185 2.120 9.515 2.735 ;
        RECT 3.190 1.970 9.515 2.120 ;
        RECT 0.115 1.950 9.515 1.970 ;
        RECT 1.870 1.800 3.520 1.950 ;
        RECT 1.870 1.780 2.040 1.800 ;
        RECT 1.565 1.550 2.040 1.780 ;
        RECT 1.565 1.130 1.805 1.550 ;
        RECT 0.615 0.770 1.805 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 1.370 2.290 1.700 3.245 ;
        RECT 2.370 2.140 3.020 3.245 ;
        RECT 3.690 2.290 4.020 3.245 ;
        RECT 4.750 2.460 6.165 2.980 ;
        RECT 6.335 2.630 6.585 3.245 ;
        RECT 6.785 2.460 7.115 2.980 ;
        RECT 7.315 2.630 7.485 3.245 ;
        RECT 7.685 2.905 9.965 3.075 ;
        RECT 7.685 2.460 8.015 2.905 ;
        RECT 4.750 2.290 8.015 2.460 ;
        RECT 8.685 2.290 9.015 2.905 ;
        RECT 9.715 1.820 9.965 2.905 ;
        RECT 5.045 1.130 9.965 1.180 ;
        RECT 0.115 0.600 0.445 1.130 ;
        RECT 1.985 0.815 3.955 1.130 ;
        RECT 4.185 1.010 9.965 1.130 ;
        RECT 4.185 0.850 6.305 1.010 ;
        RECT 4.185 0.815 4.515 0.850 ;
        RECT 1.985 0.600 2.155 0.815 ;
        RECT 5.475 0.645 5.805 0.680 ;
        RECT 0.115 0.350 2.155 0.600 ;
        RECT 2.335 0.350 5.805 0.645 ;
        RECT 5.975 0.350 6.305 0.850 ;
        RECT 6.475 0.085 6.805 0.820 ;
        RECT 6.985 0.350 7.155 1.010 ;
        RECT 7.335 0.085 7.665 0.820 ;
        RECT 7.845 0.350 8.095 1.010 ;
        RECT 8.265 0.085 8.595 0.820 ;
        RECT 8.775 0.350 9.025 1.010 ;
        RECT 9.205 0.085 9.535 0.820 ;
        RECT 9.715 0.350 9.965 1.010 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
  END
END sky130_fd_sc_hs__o2111ai_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.350 1.375 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.775 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 1.955 1.820 2.310 2.980 ;
        RECT 2.140 1.130 2.310 1.820 ;
        RECT 1.955 0.350 2.310 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.295 2.120 0.625 2.700 ;
        RECT 1.165 2.290 1.785 3.245 ;
        RECT 0.295 1.950 1.785 2.120 ;
        RECT 0.295 1.820 0.625 1.950 ;
        RECT 1.615 1.630 1.785 1.950 ;
        RECT 1.615 1.300 1.970 1.630 ;
        RECT 1.615 1.180 1.785 1.300 ;
        RECT 0.945 1.010 1.785 1.180 ;
        RECT 0.295 0.085 0.650 0.995 ;
        RECT 0.945 0.540 1.240 1.010 ;
        RECT 1.455 0.085 1.785 0.840 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__or2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.350 1.045 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.435 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 2.395 1.240 ;
        RECT 0.000 0.000 2.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 2.590 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.400 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.565600 ;
    PORT
      LAYER li1 ;
        RECT 1.555 1.820 1.835 2.150 ;
        RECT 1.555 0.350 1.795 1.820 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.400 3.415 ;
        RECT 0.105 2.490 0.435 2.860 ;
        RECT 1.035 2.660 1.365 3.245 ;
        RECT 1.955 2.660 2.285 3.245 ;
        RECT 0.105 2.320 2.295 2.490 ;
        RECT 0.105 1.820 0.435 2.320 ;
        RECT 1.215 1.180 1.385 2.320 ;
        RECT 2.125 1.630 2.295 2.320 ;
        RECT 1.965 1.300 2.295 1.630 ;
        RECT 0.620 1.010 1.385 1.180 ;
        RECT 0.110 0.085 0.440 1.000 ;
        RECT 0.620 0.450 0.870 1.010 ;
        RECT 1.045 0.085 1.375 0.825 ;
        RECT 1.970 0.085 2.300 1.130 ;
        RECT 0.000 -0.085 2.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
  END
END sky130_fd_sc_hs__or2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 2.520 1.950 3.895 2.120 ;
        RECT 2.210 1.350 2.755 1.950 ;
        RECT 3.590 1.450 3.895 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.450 3.255 1.780 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.149300 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.970 0.895 2.980 ;
        RECT 1.465 1.970 1.795 2.980 ;
        RECT 0.125 1.800 1.795 1.970 ;
        RECT 0.125 1.130 0.355 1.800 ;
        RECT 0.125 0.960 1.700 1.130 ;
        RECT 0.545 0.350 0.795 0.960 ;
        RECT 1.405 0.350 1.700 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.140 0.365 3.245 ;
        RECT 1.095 2.140 1.265 3.245 ;
        RECT 1.995 2.120 2.245 3.245 ;
        RECT 2.450 2.905 3.730 3.075 ;
        RECT 2.450 2.290 2.780 2.905 ;
        RECT 2.980 2.460 3.230 2.735 ;
        RECT 3.400 2.630 3.730 2.905 ;
        RECT 3.930 2.630 4.205 3.245 ;
        RECT 2.980 2.290 4.235 2.460 ;
        RECT 0.595 1.300 2.040 1.630 ;
        RECT 1.870 1.180 2.040 1.300 ;
        RECT 4.065 1.180 4.235 2.290 ;
        RECT 1.870 1.010 4.235 1.180 ;
        RECT 0.115 0.085 0.365 0.790 ;
        RECT 0.975 0.085 1.225 0.790 ;
        RECT 1.920 0.085 2.250 0.840 ;
        RECT 2.420 0.350 2.750 1.010 ;
        RECT 2.920 0.085 4.205 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__or2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.350 2.365 1.780 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.180 0.455 1.550 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.315 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 2.755 1.820 3.275 2.980 ;
        RECT 3.105 1.130 3.275 1.820 ;
        RECT 2.875 0.350 3.275 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 1.930 0.445 2.980 ;
        RECT 0.615 2.100 0.945 3.245 ;
        RECT 1.300 1.990 1.630 2.860 ;
        RECT 0.115 1.760 0.830 1.930 ;
        RECT 1.300 1.820 1.865 1.990 ;
        RECT 2.255 1.950 2.585 3.245 ;
        RECT 0.660 1.630 0.830 1.760 ;
        RECT 0.660 1.300 1.525 1.630 ;
        RECT 0.660 1.010 0.830 1.300 ;
        RECT 1.695 1.180 1.865 1.820 ;
        RECT 2.535 1.300 2.935 1.630 ;
        RECT 2.535 1.180 2.705 1.300 ;
        RECT 0.115 0.680 0.830 1.010 ;
        RECT 1.000 0.085 1.525 1.130 ;
        RECT 1.695 1.010 2.705 1.180 ;
        RECT 1.695 0.540 2.045 1.010 ;
        RECT 2.265 0.085 2.680 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__or2b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.350 2.365 1.780 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 1.780 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 1.140 1.900 1.240 ;
        RECT 0.010 0.245 3.355 1.140 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.787700 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.820 1.645 2.070 ;
        RECT 1.060 1.130 1.230 1.820 ;
        RECT 1.060 0.350 1.390 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.115 2.410 0.445 2.700 ;
        RECT 0.650 2.580 0.980 3.245 ;
        RECT 1.765 2.580 2.095 3.245 ;
        RECT 0.115 2.240 2.705 2.410 ;
        RECT 0.115 1.950 0.890 2.240 ;
        RECT 0.720 1.180 0.890 1.950 ;
        RECT 2.535 1.650 2.705 2.240 ;
        RECT 2.875 1.820 3.275 2.860 ;
        RECT 1.465 1.300 1.795 1.630 ;
        RECT 2.535 1.320 2.935 1.650 ;
        RECT 0.120 1.010 0.890 1.180 ;
        RECT 1.625 1.150 1.795 1.300 ;
        RECT 3.105 1.150 3.275 1.820 ;
        RECT 0.120 0.540 0.450 1.010 ;
        RECT 1.625 0.980 3.275 1.150 ;
        RECT 0.630 0.085 0.880 0.840 ;
        RECT 1.560 0.085 2.235 0.810 ;
        RECT 2.405 0.350 2.735 0.980 ;
        RECT 2.915 0.085 3.245 0.810 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__or2b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.450 3.235 1.780 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 4.905 1.120 5.235 1.790 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.140 2.335 1.240 ;
        RECT 0.005 0.245 5.570 1.140 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.104900 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.970 0.805 2.980 ;
        RECT 1.455 1.970 1.785 2.980 ;
        RECT 0.605 1.800 1.785 1.970 ;
        RECT 0.605 1.410 0.775 1.800 ;
        RECT 0.125 1.180 0.775 1.410 ;
        RECT 0.545 1.130 0.775 1.180 ;
        RECT 0.545 0.960 1.805 1.130 ;
        RECT 0.545 0.350 0.795 0.960 ;
        RECT 1.475 0.350 1.805 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.105 1.820 0.435 3.245 ;
        RECT 1.005 2.140 1.255 3.245 ;
        RECT 1.985 1.940 2.235 3.245 ;
        RECT 2.430 2.120 2.760 2.980 ;
        RECT 2.960 2.290 3.210 3.245 ;
        RECT 3.425 2.905 4.655 3.075 ;
        RECT 3.425 2.120 3.675 2.905 ;
        RECT 2.430 1.950 3.675 2.120 ;
        RECT 3.425 1.915 3.675 1.950 ;
        RECT 0.945 1.300 2.145 1.630 ;
        RECT 3.875 1.450 4.125 2.735 ;
        RECT 4.325 1.945 4.655 2.905 ;
        RECT 4.875 1.960 5.205 3.245 ;
        RECT 1.975 1.280 2.145 1.300 ;
        RECT 3.505 1.280 4.125 1.450 ;
        RECT 4.295 1.445 4.625 1.775 ;
        RECT 1.975 1.110 3.755 1.280 ;
        RECT 0.115 0.085 0.365 1.010 ;
        RECT 0.975 0.085 1.305 0.765 ;
        RECT 1.975 0.085 2.305 0.940 ;
        RECT 2.475 0.350 2.805 1.110 ;
        RECT 3.005 0.085 3.335 0.940 ;
        RECT 3.505 0.350 3.755 1.110 ;
        RECT 3.935 0.085 4.265 1.030 ;
        RECT 4.435 0.950 4.625 1.445 ;
        RECT 5.405 0.950 5.655 2.980 ;
        RECT 4.435 0.350 5.655 0.950 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__or2b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.350 1.815 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.350 1.315 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.570 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 2.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.925 1.050 2.870 1.240 ;
        RECT 0.005 0.245 2.870 1.050 ;
        RECT 0.000 0.000 2.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 2.880 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.820 2.795 2.980 ;
        RECT 2.625 1.130 2.795 1.820 ;
        RECT 2.430 0.350 2.795 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.115 2.120 0.445 2.860 ;
        RECT 1.555 2.290 2.315 3.245 ;
        RECT 0.115 1.950 2.260 2.120 ;
        RECT 2.090 1.630 2.260 1.950 ;
        RECT 2.090 1.300 2.455 1.630 ;
        RECT 2.090 1.180 2.260 1.300 ;
        RECT 0.115 1.010 2.260 1.180 ;
        RECT 0.115 0.350 0.365 1.010 ;
        RECT 0.545 0.085 0.875 0.810 ;
        RECT 1.045 0.455 1.760 1.010 ;
        RECT 1.930 0.085 2.260 0.810 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
  END
END sky130_fd_sc_hs__or3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.180 1.905 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.130 1.335 2.890 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.120 0.835 1.790 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.910 1.140 3.355 1.240 ;
        RECT 0.005 0.245 3.355 1.140 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.970 2.665 2.980 ;
        RECT 2.335 1.800 3.235 1.970 ;
        RECT 3.005 1.130 3.235 1.800 ;
        RECT 2.415 0.960 3.235 1.130 ;
        RECT 2.415 0.350 2.745 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.285 2.130 0.615 2.980 ;
        RECT 0.095 1.960 0.615 2.130 ;
        RECT 0.095 0.950 0.265 1.960 ;
        RECT 1.725 1.940 2.055 3.245 ;
        RECT 2.835 2.140 3.165 3.245 ;
        RECT 2.075 1.300 2.815 1.630 ;
        RECT 2.075 0.960 2.245 1.300 ;
        RECT 1.200 0.950 2.245 0.960 ;
        RECT 0.095 0.790 2.245 0.950 ;
        RECT 0.095 0.780 1.530 0.790 ;
        RECT 0.095 0.350 0.445 0.780 ;
        RECT 0.615 0.085 1.030 0.600 ;
        RECT 1.200 0.350 1.530 0.780 ;
        RECT 1.700 0.085 2.245 0.600 ;
        RECT 2.915 0.085 3.245 0.790 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__or3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.280 0.435 1.630 ;
        RECT 2.755 1.280 3.055 1.550 ;
        RECT 0.105 1.110 3.055 1.280 ;
        RECT 0.105 0.280 0.435 1.110 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.450 2.545 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.270 1.380 0.940 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.440 0.245 5.275 1.240 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.090100 ;
    PORT
      LAYER li1 ;
        RECT 3.565 1.970 3.735 2.980 ;
        RECT 4.385 1.970 4.715 2.980 ;
        RECT 3.565 1.800 5.155 1.970 ;
        RECT 4.925 1.130 5.155 1.800 ;
        RECT 3.565 0.960 5.155 1.130 ;
        RECT 3.565 0.350 3.735 0.960 ;
        RECT 4.405 0.350 4.655 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.115 1.920 0.365 3.245 ;
        RECT 0.565 2.540 0.815 2.960 ;
        RECT 1.015 2.710 2.330 2.960 ;
        RECT 2.500 2.540 2.830 2.960 ;
        RECT 0.565 2.370 2.830 2.540 ;
        RECT 0.565 1.950 0.815 2.370 ;
        RECT 2.500 2.290 2.830 2.370 ;
        RECT 3.035 2.290 3.365 3.245 ;
        RECT 1.495 2.120 1.825 2.200 ;
        RECT 3.935 2.140 4.185 3.245 ;
        RECT 4.915 2.140 5.165 3.245 ;
        RECT 1.495 1.950 3.395 2.120 ;
        RECT 3.225 1.630 3.395 1.950 ;
        RECT 3.225 1.300 4.685 1.630 ;
        RECT 3.225 0.940 3.395 1.300 ;
        RECT 1.550 0.770 3.395 0.940 ;
        RECT 1.550 0.350 1.880 0.770 ;
        RECT 2.050 0.085 2.380 0.600 ;
        RECT 2.550 0.350 2.880 0.770 ;
        RECT 3.050 0.085 3.380 0.600 ;
        RECT 3.915 0.085 4.165 0.790 ;
        RECT 4.835 0.085 5.165 0.790 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__or3_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.300 2.845 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 1.915 1.190 2.275 2.890 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.110 0.605 1.780 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.890 1.050 3.835 1.240 ;
        RECT 0.005 0.245 3.835 1.050 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.250 1.820 3.755 2.980 ;
        RECT 3.585 1.130 3.755 1.820 ;
        RECT 3.395 0.350 3.755 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 2.100 0.445 3.245 ;
        RECT 0.615 2.100 0.945 2.980 ;
        RECT 0.775 1.880 0.945 2.100 ;
        RECT 0.775 1.210 1.205 1.880 ;
        RECT 0.775 0.940 0.945 1.210 ;
        RECT 1.375 1.020 1.705 2.975 ;
        RECT 2.750 1.950 3.080 3.245 ;
        RECT 3.055 1.300 3.415 1.630 ;
        RECT 3.055 1.020 3.225 1.300 ;
        RECT 0.115 0.085 0.445 0.940 ;
        RECT 0.615 0.350 0.945 0.940 ;
        RECT 1.175 0.850 3.225 1.020 ;
        RECT 1.175 0.350 1.505 0.850 ;
        RECT 1.675 0.085 2.005 0.680 ;
        RECT 2.175 0.350 2.505 0.850 ;
        RECT 2.675 0.085 3.225 0.680 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__or3b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.350 2.305 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.350 2.845 1.780 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.300 0.435 1.780 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.075 0.245 3.790 1.240 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.820 1.795 2.150 ;
        RECT 1.065 1.130 1.235 1.820 ;
        RECT 1.065 0.960 1.455 1.130 ;
        RECT 1.125 0.350 1.455 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.115 2.490 0.445 2.700 ;
        RECT 0.650 2.660 0.980 3.245 ;
        RECT 1.635 2.660 2.070 3.245 ;
        RECT 0.115 2.320 2.645 2.490 ;
        RECT 0.115 1.950 0.775 2.320 ;
        RECT 2.475 2.120 2.645 2.320 ;
        RECT 3.235 2.290 3.755 2.860 ;
        RECT 2.475 1.950 3.415 2.120 ;
        RECT 0.605 1.130 0.775 1.950 ;
        RECT 1.405 1.300 1.795 1.630 ;
        RECT 3.085 1.350 3.415 1.950 ;
        RECT 0.185 0.960 0.775 1.130 ;
        RECT 1.625 1.180 1.795 1.300 ;
        RECT 3.585 1.180 3.755 2.290 ;
        RECT 1.625 1.010 3.755 1.180 ;
        RECT 0.185 0.540 0.605 0.960 ;
        RECT 0.775 0.085 0.945 0.790 ;
        RECT 1.625 0.085 2.135 0.780 ;
        RECT 2.350 0.450 2.680 1.010 ;
        RECT 2.850 0.085 3.180 0.840 ;
        RECT 3.350 0.450 3.755 1.010 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__or3b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 0.800 1.320 1.130 1.760 ;
        RECT 3.285 1.380 3.545 1.550 ;
        RECT 3.005 1.320 3.545 1.380 ;
        RECT 0.800 1.150 3.545 1.320 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 1.340 1.550 3.075 1.800 ;
        RECT 1.340 1.490 1.670 1.550 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 0.775 0.640 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 1.240 1.520 1.450 ;
        RECT 0.025 0.245 5.755 1.240 ;
        RECT 0.000 0.000 5.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.760 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.104900 ;
    PORT
      LAYER li1 ;
        RECT 4.055 1.970 4.225 2.980 ;
        RECT 4.875 1.970 5.205 2.980 ;
        RECT 4.055 1.800 5.635 1.970 ;
        RECT 5.405 1.130 5.635 1.800 ;
        RECT 4.055 0.960 5.635 1.130 ;
        RECT 4.055 0.350 4.225 0.960 ;
        RECT 4.885 0.350 5.135 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.760 3.415 ;
        RECT 0.110 1.340 0.360 2.980 ;
        RECT 0.560 1.940 0.890 3.245 ;
        RECT 1.070 2.530 1.400 2.980 ;
        RECT 1.580 2.700 2.835 2.980 ;
        RECT 3.005 2.530 3.335 2.980 ;
        RECT 1.070 2.360 3.335 2.530 ;
        RECT 1.070 1.970 1.400 2.360 ;
        RECT 3.005 2.310 3.335 2.360 ;
        RECT 3.505 2.310 3.835 3.245 ;
        RECT 2.030 2.140 2.385 2.190 ;
        RECT 4.425 2.140 4.675 3.245 ;
        RECT 5.405 2.140 5.655 3.245 ;
        RECT 2.030 1.970 3.885 2.140 ;
        RECT 3.715 1.630 3.885 1.970 ;
        RECT 0.110 0.980 0.465 1.340 ;
        RECT 3.715 1.300 5.175 1.630 ;
        RECT 3.715 0.980 3.885 1.300 ;
        RECT 0.110 0.810 1.910 0.980 ;
        RECT 0.945 0.085 1.410 0.640 ;
        RECT 1.580 0.310 1.910 0.810 ;
        RECT 2.080 0.810 3.885 0.980 ;
        RECT 2.080 0.350 2.410 0.810 ;
        RECT 2.580 0.085 2.910 0.640 ;
        RECT 3.090 0.350 3.340 0.810 ;
        RECT 3.510 0.085 3.850 0.600 ;
        RECT 4.405 0.085 4.655 0.790 ;
        RECT 5.315 0.085 5.645 0.790 ;
        RECT 0.000 -0.085 5.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
  END
END sky130_fd_sc_hs__or3b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.390 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.420 1.820 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 0.920 1.420 1.295 1.780 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.420 0.650 1.780 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 3.320 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 2.900 1.820 3.275 2.980 ;
        RECT 3.105 1.130 3.275 1.820 ;
        RECT 2.960 0.350 3.275 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.200 2.120 0.530 2.980 ;
        RECT 2.150 2.290 2.565 3.245 ;
        RECT 0.200 1.950 2.730 2.120 ;
        RECT 2.560 1.630 2.730 1.950 ;
        RECT 2.560 1.300 2.935 1.630 ;
        RECT 2.560 1.180 2.730 1.300 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 0.615 1.010 2.730 1.180 ;
        RECT 0.615 0.540 0.945 1.010 ;
        RECT 1.125 0.085 1.600 0.840 ;
        RECT 1.860 0.540 2.190 1.010 ;
        RECT 2.450 0.085 2.780 0.840 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__or4_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.350 2.455 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.350 1.875 2.890 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.165 1.335 2.890 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.180 0.835 1.770 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.460 1.140 3.835 1.240 ;
        RECT 0.005 0.245 3.835 1.140 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 2.860 1.970 3.190 2.980 ;
        RECT 2.860 1.800 3.715 1.970 ;
        RECT 3.485 1.130 3.715 1.800 ;
        RECT 2.965 0.960 3.715 1.130 ;
        RECT 2.965 0.350 3.215 0.960 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.405 2.110 0.735 2.980 ;
        RECT 0.085 1.940 0.735 2.110 ;
        RECT 2.360 1.950 2.690 3.245 ;
        RECT 3.360 2.140 3.690 3.245 ;
        RECT 0.085 0.995 0.255 1.940 ;
        RECT 2.625 1.300 3.040 1.630 ;
        RECT 2.625 1.180 2.795 1.300 ;
        RECT 1.860 1.010 2.795 1.180 ;
        RECT 1.860 0.995 2.190 1.010 ;
        RECT 0.085 0.825 2.190 0.995 ;
        RECT 0.115 0.085 0.510 0.655 ;
        RECT 0.690 0.350 1.020 0.825 ;
        RECT 1.200 0.085 1.680 0.655 ;
        RECT 1.860 0.350 2.190 0.825 ;
        RECT 2.360 0.085 2.795 0.825 ;
        RECT 3.395 0.085 3.725 0.775 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__or4_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.470 3.735 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.410 3.235 1.550 ;
        RECT 2.525 1.300 3.235 1.410 ;
        RECT 4.065 1.300 4.395 1.550 ;
        RECT 2.525 1.130 4.395 1.300 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.770 6.285 1.780 ;
        RECT 4.605 1.365 6.285 1.770 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 6.285 0.255 6.615 0.855 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 6.720 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.790 5.675 1.240 ;
        RECT 0.005 0.245 6.225 0.790 ;
        RECT 0.000 0.000 6.720 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 6.910 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 6.720 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.326900 ;
    PORT
      LAYER li1 ;
        RECT 0.615 2.150 0.845 2.980 ;
        RECT 1.515 2.150 1.745 2.980 ;
        RECT 0.125 1.820 2.275 2.150 ;
        RECT 0.125 1.300 0.945 1.820 ;
        RECT 0.615 1.150 0.945 1.300 ;
        RECT 0.615 0.980 1.945 1.150 ;
        RECT 0.615 0.350 0.945 0.980 ;
        RECT 1.615 0.350 1.945 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 6.720 3.415 ;
        RECT 0.115 2.320 0.445 3.245 ;
        RECT 1.015 2.320 1.345 3.245 ;
        RECT 1.915 2.320 2.245 3.245 ;
        RECT 2.475 2.190 2.755 2.980 ;
        RECT 2.925 2.560 3.205 2.980 ;
        RECT 3.375 2.730 3.705 3.245 ;
        RECT 3.895 2.560 4.175 2.980 ;
        RECT 2.925 2.360 4.175 2.560 ;
        RECT 3.825 2.310 4.175 2.360 ;
        RECT 4.345 2.530 4.675 2.980 ;
        RECT 4.845 2.700 6.075 2.980 ;
        RECT 6.245 2.530 6.575 2.980 ;
        RECT 4.345 2.360 6.575 2.530 ;
        RECT 2.475 2.140 2.805 2.190 ;
        RECT 4.345 2.140 4.675 2.360 ;
        RECT 6.245 2.290 6.575 2.360 ;
        RECT 2.475 1.970 4.675 2.140 ;
        RECT 2.475 1.940 2.805 1.970 ;
        RECT 4.345 1.940 4.675 1.970 ;
        RECT 5.295 2.120 5.625 2.190 ;
        RECT 5.295 1.950 6.635 2.120 ;
        RECT 1.315 1.320 2.325 1.650 ;
        RECT 0.115 0.085 0.445 1.130 ;
        RECT 2.155 0.960 2.325 1.320 ;
        RECT 6.465 1.195 6.635 1.950 ;
        RECT 4.770 1.025 6.635 1.195 ;
        RECT 4.770 0.960 5.100 1.025 ;
        RECT 1.115 0.085 1.445 0.810 ;
        RECT 2.155 0.790 5.100 0.960 ;
        RECT 2.380 0.085 2.740 0.620 ;
        RECT 2.920 0.350 3.250 0.790 ;
        RECT 3.430 0.085 4.590 0.620 ;
        RECT 4.770 0.350 5.100 0.790 ;
        RECT 5.270 0.085 6.115 0.680 ;
        RECT 0.000 -0.085 6.720 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
  END
END sky130_fd_sc_hs__or4_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.995 1.350 3.325 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.455 1.180 2.785 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.045 2.275 1.780 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.450 0.570 1.780 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.330 1.050 4.275 1.240 ;
        RECT 0.005 0.245 4.275 1.050 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 3.835 1.820 4.235 2.980 ;
        RECT 4.065 1.130 4.235 1.820 ;
        RECT 3.835 0.350 4.235 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.120 2.120 0.450 2.980 ;
        RECT 0.620 2.290 0.950 3.245 ;
        RECT 1.315 2.120 1.645 2.860 ;
        RECT 3.335 2.290 3.665 3.245 ;
        RECT 0.120 1.950 0.980 2.120 ;
        RECT 0.810 1.910 0.980 1.950 ;
        RECT 1.315 1.950 3.665 2.120 ;
        RECT 0.810 1.580 1.140 1.910 ;
        RECT 0.810 1.280 0.980 1.580 ;
        RECT 0.115 1.110 0.980 1.280 ;
        RECT 0.115 0.350 0.445 1.110 ;
        RECT 0.615 0.085 0.945 0.940 ;
        RECT 1.315 0.875 1.645 1.950 ;
        RECT 3.495 1.630 3.665 1.950 ;
        RECT 3.495 1.300 3.895 1.630 ;
        RECT 3.495 1.180 3.665 1.300 ;
        RECT 2.955 1.010 3.665 1.180 ;
        RECT 2.955 0.940 3.125 1.010 ;
        RECT 1.115 0.545 2.090 0.875 ;
        RECT 2.260 0.085 2.590 0.875 ;
        RECT 2.760 0.350 3.125 0.940 ;
        RECT 3.295 0.085 3.625 0.840 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__or4b_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.350 2.275 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.470 2.815 2.150 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.470 3.355 2.520 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 1.780 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.245 4.315 1.240 ;
        RECT 0.000 0.000 4.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.320 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.820 1.430 2.150 ;
        RECT 1.060 1.130 1.230 1.820 ;
        RECT 1.060 0.350 1.405 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.115 2.490 0.445 2.700 ;
        RECT 0.650 2.660 0.980 3.245 ;
        RECT 1.550 2.730 2.125 3.245 ;
        RECT 2.295 2.690 3.695 2.860 ;
        RECT 2.295 2.490 2.465 2.690 ;
        RECT 0.115 2.320 2.465 2.490 ;
        RECT 0.115 1.950 0.890 2.320 ;
        RECT 0.720 1.180 0.890 1.950 ;
        RECT 3.525 1.770 3.695 2.690 ;
        RECT 3.865 1.940 4.235 2.980 ;
        RECT 1.400 1.300 1.745 1.630 ;
        RECT 3.525 1.440 3.895 1.770 ;
        RECT 0.130 1.010 0.890 1.180 ;
        RECT 1.575 1.130 1.745 1.300 ;
        RECT 4.065 1.270 4.235 1.940 ;
        RECT 3.375 1.130 4.235 1.270 ;
        RECT 1.575 1.100 4.235 1.130 ;
        RECT 0.130 0.540 0.460 1.010 ;
        RECT 1.575 0.960 3.705 1.100 ;
        RECT 0.640 0.085 0.890 0.840 ;
        RECT 1.575 0.085 1.995 0.780 ;
        RECT 2.175 0.450 2.505 0.960 ;
        RECT 2.685 0.085 3.205 0.780 ;
        RECT 3.375 0.450 3.705 0.960 ;
        RECT 3.875 0.085 4.205 0.930 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
  END
END sky130_fd_sc_hs__or4b_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.450 1.335 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.280 0.835 1.550 ;
        RECT 1.705 1.280 2.035 1.550 ;
        RECT 0.125 1.110 2.035 1.280 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 2.495 1.365 2.785 1.410 ;
        RECT 3.935 1.365 4.225 1.410 ;
        RECT 2.495 1.225 4.225 1.365 ;
        RECT 2.495 1.180 2.785 1.225 ;
        RECT 3.935 1.180 4.225 1.225 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.180 4.815 1.550 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.200 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.780 3.380 1.240 ;
        RECT 4.240 0.780 7.195 1.240 ;
        RECT 0.005 0.245 7.195 0.780 ;
        RECT 0.000 0.000 7.200 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.390 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.200 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.178900 ;
    PORT
      LAYER li1 ;
        RECT 5.410 2.150 5.690 2.980 ;
        RECT 6.360 2.150 6.590 2.980 ;
        RECT 5.410 1.820 7.075 2.150 ;
        RECT 6.365 1.470 6.655 1.820 ;
        RECT 6.325 1.300 6.655 1.470 ;
        RECT 6.325 1.150 6.575 1.300 ;
        RECT 5.325 0.980 6.575 1.150 ;
        RECT 5.325 0.350 5.655 0.980 ;
        RECT 6.325 0.350 6.575 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.115 2.120 0.445 2.980 ;
        RECT 0.645 2.460 0.815 2.980 ;
        RECT 1.015 2.630 1.345 3.245 ;
        RECT 1.515 2.460 1.845 2.980 ;
        RECT 0.645 2.290 1.845 2.460 ;
        RECT 2.015 2.530 2.345 2.980 ;
        RECT 2.515 2.700 3.745 2.980 ;
        RECT 3.945 2.530 4.195 2.980 ;
        RECT 2.015 2.360 4.195 2.530 ;
        RECT 2.015 2.120 2.345 2.360 ;
        RECT 0.115 1.950 2.345 2.120 ;
        RECT 2.895 2.020 3.295 2.190 ;
        RECT 3.945 2.060 4.195 2.360 ;
        RECT 0.115 1.940 0.445 1.950 ;
        RECT 2.245 1.180 2.725 1.780 ;
        RECT 2.895 1.130 3.065 2.020 ;
        RECT 4.425 1.890 4.755 2.860 ;
        RECT 3.465 1.800 4.755 1.890 ;
        RECT 4.960 1.820 5.210 3.245 ;
        RECT 5.860 2.320 6.190 3.245 ;
        RECT 6.760 2.320 7.090 3.245 ;
        RECT 3.235 1.720 4.755 1.800 ;
        RECT 3.235 1.470 3.635 1.720 ;
        RECT 3.865 1.180 4.195 1.510 ;
        RECT 4.985 1.320 6.155 1.650 ;
        RECT 2.895 1.010 3.270 1.130 ;
        RECT 4.985 1.010 5.155 1.320 ;
        RECT 2.895 0.940 5.155 1.010 ;
        RECT 0.115 0.840 5.155 0.940 ;
        RECT 0.115 0.770 3.270 0.840 ;
        RECT 0.115 0.350 0.445 0.770 ;
        RECT 0.615 0.085 0.945 0.600 ;
        RECT 1.115 0.350 2.200 0.770 ;
        RECT 2.370 0.085 2.725 0.600 ;
        RECT 2.895 0.350 3.270 0.770 ;
        RECT 3.440 0.340 4.565 0.670 ;
        RECT 4.825 0.085 5.155 0.670 ;
        RECT 5.825 0.085 6.155 0.810 ;
        RECT 6.755 0.085 7.085 1.130 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 2.555 1.210 2.725 1.380 ;
        RECT 3.995 1.210 4.165 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
  END
END sky130_fd_sc_hs__or4b_4

#--------EOF---------

MACRO sky130_fd_sc_hs__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 3.835 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.232500 ;
    PORT
      LAYER li1 ;
        RECT 2.965 1.350 3.295 2.890 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.300 0.455 1.780 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.050 1.315 1.720 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.840 1.050 4.785 1.240 ;
        RECT 0.030 0.245 4.785 1.050 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 4.240 1.820 4.715 2.980 ;
        RECT 4.545 1.130 4.715 1.820 ;
        RECT 4.345 0.350 4.715 1.130 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 2.480 0.445 2.980 ;
        RECT 0.615 2.650 0.945 3.245 ;
        RECT 1.115 2.905 2.755 3.075 ;
        RECT 1.115 2.480 1.285 2.905 ;
        RECT 0.115 2.310 1.285 2.480 ;
        RECT 0.115 2.100 0.795 2.310 ;
        RECT 0.625 1.130 0.795 2.100 ;
        RECT 1.150 1.890 1.655 2.140 ;
        RECT 0.140 0.960 0.795 1.130 ;
        RECT 1.485 1.700 1.655 1.890 ;
        RECT 1.845 1.870 2.245 2.735 ;
        RECT 1.485 1.030 1.905 1.700 ;
        RECT 0.140 0.350 0.470 0.960 ;
        RECT 1.485 0.880 1.655 1.030 ;
        RECT 0.640 0.085 0.970 0.790 ;
        RECT 1.140 0.350 1.655 0.880 ;
        RECT 2.075 1.020 2.245 1.870 ;
        RECT 2.425 1.190 2.755 2.905 ;
        RECT 3.740 1.950 4.070 3.245 ;
        RECT 4.005 1.300 4.375 1.630 ;
        RECT 4.005 1.180 4.175 1.300 ;
        RECT 3.310 1.020 4.175 1.180 ;
        RECT 2.075 1.010 4.175 1.020 ;
        RECT 2.075 0.850 3.640 1.010 ;
        RECT 1.825 0.085 2.075 0.680 ;
        RECT 2.245 0.350 2.575 0.850 ;
        RECT 2.745 0.085 3.140 0.680 ;
        RECT 3.310 0.350 3.640 0.850 ;
        RECT 3.810 0.085 4.140 0.840 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__or4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hs__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.470 3.925 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.570 3.715 0.670 ;
        RECT 3.150 0.255 3.715 0.570 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 1.300 4.695 1.780 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.350 0.550 1.780 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.200 1.370 4.250 1.450 ;
        RECT 0.010 1.135 4.250 1.370 ;
        RECT 0.010 0.245 4.795 1.135 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.850 1.390 2.100 ;
        RECT 1.060 1.180 1.230 1.850 ;
        RECT 1.060 0.440 1.315 1.180 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.105 2.440 0.435 2.980 ;
        RECT 0.605 2.610 0.935 3.245 ;
        RECT 1.510 2.610 1.840 3.245 ;
        RECT 2.050 2.780 2.380 2.980 ;
        RECT 2.050 2.610 2.605 2.780 ;
        RECT 0.105 2.270 2.265 2.440 ;
        RECT 0.105 2.100 0.890 2.270 ;
        RECT 0.720 1.180 0.890 2.100 ;
        RECT 1.400 1.350 1.730 1.680 ;
        RECT 1.970 1.470 2.265 2.270 ;
        RECT 0.120 1.010 0.890 1.180 ;
        RECT 1.560 1.300 1.730 1.350 ;
        RECT 2.435 1.300 2.605 2.610 ;
        RECT 3.820 2.310 4.150 3.245 ;
        RECT 4.360 2.140 4.690 2.820 ;
        RECT 2.775 1.970 4.690 2.140 ;
        RECT 2.775 1.470 3.070 1.970 ;
        RECT 4.095 1.950 4.690 1.970 ;
        RECT 1.560 1.130 3.735 1.300 ;
        RECT 0.120 0.670 0.450 1.010 ;
        RECT 0.630 0.085 0.880 0.840 ;
        RECT 1.575 0.085 2.035 0.910 ;
        RECT 2.310 0.580 2.640 1.130 ;
        RECT 2.810 0.740 3.195 0.960 ;
        RECT 3.405 0.840 3.735 1.130 ;
        RECT 4.095 1.130 4.265 1.950 ;
        RECT 4.095 0.960 4.685 1.130 ;
        RECT 2.810 0.085 2.980 0.740 ;
        RECT 3.925 0.085 4.255 0.790 ;
        RECT 4.435 0.435 4.685 0.960 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__or4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hs__or4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 7.525 1.180 8.535 1.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.450 7.075 1.780 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.375 1.350 3.715 1.780 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.350 0.835 1.780 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.245 8.420 1.240 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.677500 ;
    PORT
      LAYER li1 ;
        RECT 1.085 2.050 2.525 2.220 ;
        RECT 1.085 1.180 1.450 2.050 ;
        RECT 1.120 0.750 1.450 1.180 ;
        RECT 1.120 0.580 2.775 0.750 ;
        RECT 1.120 0.350 1.450 0.580 ;
        RECT 2.140 0.420 2.775 0.580 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.085 2.560 0.445 2.860 ;
        RECT 0.650 2.730 0.995 3.245 ;
        RECT 1.565 2.730 1.990 3.245 ;
        RECT 2.840 2.730 3.170 3.245 ;
        RECT 4.835 2.980 6.115 3.075 ;
        RECT 3.935 2.905 6.115 2.980 ;
        RECT 3.935 2.630 5.165 2.905 ;
        RECT 0.085 2.390 2.865 2.560 ;
        RECT 0.085 1.950 0.445 2.390 ;
        RECT 0.085 1.130 0.255 1.950 ;
        RECT 2.695 1.880 2.865 2.390 ;
        RECT 1.620 1.710 2.865 1.880 ;
        RECT 3.035 2.290 4.715 2.460 ;
        RECT 0.085 0.450 0.445 1.130 ;
        RECT 0.615 0.085 0.915 1.130 ;
        RECT 1.620 1.090 1.790 1.710 ;
        RECT 3.035 1.540 3.205 2.290 ;
        RECT 3.375 1.950 4.055 2.120 ;
        RECT 1.960 1.260 3.205 1.540 ;
        RECT 3.885 1.590 4.055 1.950 ;
        RECT 4.385 1.930 4.715 2.290 ;
        RECT 5.335 2.270 5.665 2.735 ;
        RECT 5.865 2.440 6.115 2.905 ;
        RECT 6.345 2.905 7.575 3.075 ;
        RECT 6.345 2.440 6.675 2.905 ;
        RECT 6.875 2.270 7.045 2.735 ;
        RECT 5.335 2.100 7.045 2.270 ;
        RECT 6.575 1.950 7.045 2.100 ;
        RECT 7.245 2.240 7.575 2.905 ;
        RECT 7.745 2.410 8.075 3.245 ;
        RECT 8.250 2.240 8.525 2.990 ;
        RECT 7.245 1.950 8.525 2.240 ;
        RECT 8.195 1.940 8.525 1.950 ;
        RECT 4.385 1.760 6.145 1.930 ;
        RECT 3.885 1.420 5.805 1.590 ;
        RECT 4.445 1.260 5.805 1.420 ;
        RECT 5.975 1.260 6.145 1.760 ;
        RECT 3.945 1.090 4.275 1.250 ;
        RECT 1.620 0.920 4.275 1.090 ;
        RECT 4.445 0.750 4.615 1.260 ;
        RECT 5.975 1.090 7.355 1.260 ;
        RECT 1.630 0.085 1.960 0.410 ;
        RECT 2.945 0.085 3.275 0.750 ;
        RECT 3.455 0.580 4.615 0.750 ;
        RECT 3.455 0.450 3.785 0.580 ;
        RECT 4.015 0.085 4.605 0.410 ;
        RECT 4.785 0.350 6.280 1.090 ;
        RECT 6.450 0.085 6.780 0.920 ;
        RECT 7.025 0.350 7.355 1.090 ;
        RECT 7.640 0.085 8.310 0.985 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__or4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfbbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.470 1.350 3.800 1.780 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.480 1.815 1.810 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 14.075 1.190 14.380 1.550 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.205 0.550 1.875 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.205 1.315 1.875 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER met1 ;
        RECT 8.255 2.105 8.545 2.150 ;
        RECT 11.615 2.105 11.905 2.150 ;
        RECT 8.255 1.965 11.905 2.105 ;
        RECT 8.255 1.920 8.545 1.965 ;
        RECT 11.615 1.920 11.905 1.965 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 16.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.180 1.145 4.900 1.280 ;
        RECT 7.040 1.240 10.690 1.275 ;
        RECT 7.040 1.145 16.775 1.240 ;
        RECT 0.030 0.245 16.775 1.145 ;
        RECT 0.000 0.000 16.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.990 3.520 ;
        RECT 13.420 1.550 15.300 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 16.800 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 16.355 1.820 16.715 2.980 ;
        RECT 16.545 1.050 16.715 1.820 ;
        RECT 16.335 0.350 16.715 1.050 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 14.890 1.820 15.275 2.980 ;
        RECT 15.105 1.130 15.275 1.820 ;
        RECT 14.915 0.350 15.275 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 16.800 3.415 ;
        RECT 0.115 2.215 0.395 2.980 ;
        RECT 0.565 2.385 0.895 3.245 ;
        RECT 1.065 2.905 2.245 3.075 ;
        RECT 1.065 2.215 1.235 2.905 ;
        RECT 1.465 2.300 1.715 2.735 ;
        RECT 1.915 2.320 2.245 2.905 ;
        RECT 2.470 2.300 2.720 3.245 ;
        RECT 2.890 2.300 3.250 2.980 ;
        RECT 0.115 2.045 1.235 2.215 ;
        RECT 1.545 2.150 1.715 2.300 ;
        RECT 1.545 1.980 2.155 2.150 ;
        RECT 1.985 1.310 2.155 1.980 ;
        RECT 2.890 1.810 3.060 2.300 ;
        RECT 3.480 2.120 3.730 2.980 ;
        RECT 3.930 2.290 4.180 3.245 ;
        RECT 3.480 1.950 4.140 2.120 ;
        RECT 2.510 1.480 3.060 1.810 ;
        RECT 1.485 1.140 2.560 1.310 ;
        RECT 1.485 1.035 1.655 1.140 ;
        RECT 0.140 0.085 0.470 1.035 ;
        RECT 0.960 0.865 1.655 1.035 ;
        RECT 0.960 0.575 1.290 0.865 ;
        RECT 1.890 0.085 2.220 0.970 ;
        RECT 2.390 0.425 2.560 1.140 ;
        RECT 2.730 0.595 3.060 1.480 ;
        RECT 3.970 1.670 4.140 1.950 ;
        RECT 4.380 1.840 4.780 2.980 ;
        RECT 5.020 2.465 5.270 3.245 ;
        RECT 5.440 2.905 7.505 3.075 ;
        RECT 5.440 2.295 5.610 2.905 ;
        RECT 6.925 2.820 7.505 2.905 ;
        RECT 4.950 2.125 5.610 2.295 ;
        RECT 5.865 2.245 6.195 2.735 ;
        RECT 6.365 2.480 6.695 2.735 ;
        RECT 6.925 2.650 7.930 2.820 ;
        RECT 8.125 2.650 8.295 3.245 ;
        RECT 7.760 2.480 7.930 2.650 ;
        RECT 8.495 2.480 8.830 2.980 ;
        RECT 6.365 2.310 7.590 2.480 ;
        RECT 6.025 2.140 6.195 2.245 ;
        RECT 4.950 1.965 5.215 2.125 ;
        RECT 6.025 1.970 7.250 2.140 ;
        RECT 4.610 1.720 4.780 1.840 ;
        RECT 5.405 1.800 5.755 1.905 ;
        RECT 5.405 1.720 6.710 1.800 ;
        RECT 3.970 1.340 4.440 1.670 ;
        RECT 4.610 1.550 6.710 1.720 ;
        RECT 3.970 1.170 4.140 1.340 ;
        RECT 4.610 1.170 4.790 1.550 ;
        RECT 6.380 1.470 6.710 1.550 ;
        RECT 3.290 0.920 4.140 1.170 ;
        RECT 4.310 0.920 4.790 1.170 ;
        RECT 4.960 1.205 5.970 1.375 ;
        RECT 6.920 1.300 7.250 1.970 ;
        RECT 4.960 0.750 5.130 1.205 ;
        RECT 3.230 0.580 5.130 0.750 ;
        RECT 3.230 0.425 3.400 0.580 ;
        RECT 2.390 0.255 3.400 0.425 ;
        RECT 3.800 0.085 4.130 0.410 ;
        RECT 5.300 0.085 5.630 1.035 ;
        RECT 5.800 0.425 5.970 1.205 ;
        RECT 6.170 1.130 7.250 1.300 ;
        RECT 6.170 0.595 6.420 1.130 ;
        RECT 7.420 0.960 7.590 2.310 ;
        RECT 6.595 0.790 7.590 0.960 ;
        RECT 7.760 2.310 8.830 2.480 ;
        RECT 9.050 2.470 9.380 3.245 ;
        RECT 7.760 1.080 7.930 2.310 ;
        RECT 8.660 2.300 8.830 2.310 ;
        RECT 8.285 1.960 8.490 2.140 ;
        RECT 8.660 2.130 9.530 2.300 ;
        RECT 8.285 1.790 8.990 1.960 ;
        RECT 8.660 1.630 8.990 1.790 ;
        RECT 9.200 1.630 9.530 2.130 ;
        RECT 9.890 2.280 10.220 2.980 ;
        RECT 10.900 2.970 11.230 3.245 ;
        RECT 11.460 2.800 11.790 2.980 ;
        RECT 11.995 2.970 12.325 3.245 ;
        RECT 12.950 2.800 13.280 2.980 ;
        RECT 10.665 2.630 13.280 2.800 ;
        RECT 9.890 2.110 10.410 2.280 ;
        RECT 8.100 1.460 8.430 1.620 ;
        RECT 9.725 1.555 10.070 1.940 ;
        RECT 10.240 1.895 10.410 2.110 ;
        RECT 10.665 2.065 10.995 2.630 ;
        RECT 11.170 2.290 12.780 2.460 ;
        RECT 11.170 1.895 11.340 2.290 ;
        RECT 10.240 1.725 11.340 1.895 ;
        RECT 8.100 1.290 9.555 1.460 ;
        RECT 6.595 0.425 6.925 0.790 ;
        RECT 5.800 0.255 6.925 0.425 ;
        RECT 7.150 0.425 7.480 0.620 ;
        RECT 7.760 0.595 8.090 1.080 ;
        RECT 8.260 0.425 8.590 1.080 ;
        RECT 7.150 0.255 8.590 0.425 ;
        RECT 8.795 0.085 9.125 1.080 ;
        RECT 9.385 0.535 9.555 1.290 ;
        RECT 9.725 1.260 11.000 1.555 ;
        RECT 11.170 1.090 11.340 1.725 ;
        RECT 11.630 1.470 11.960 2.120 ;
        RECT 12.610 1.890 12.780 2.290 ;
        RECT 12.950 2.380 13.280 2.630 ;
        RECT 14.000 2.550 14.690 3.245 ;
        RECT 12.950 2.210 14.720 2.380 ;
        RECT 12.950 2.060 13.280 2.210 ;
        RECT 12.610 1.720 13.440 1.890 ;
        RECT 12.200 1.300 12.530 1.550 ;
        RECT 12.770 1.470 13.440 1.720 ;
        RECT 13.610 1.790 14.130 2.040 ;
        RECT 13.610 1.300 13.780 1.790 ;
        RECT 14.550 1.630 14.720 2.210 ;
        RECT 14.550 1.300 14.935 1.630 ;
        RECT 15.450 1.550 15.700 2.780 ;
        RECT 15.905 1.900 16.155 3.245 ;
        RECT 9.745 0.920 11.340 1.090 ;
        RECT 11.510 1.130 13.905 1.300 ;
        RECT 9.745 0.705 10.580 0.920 ;
        RECT 11.510 0.750 11.680 1.130 ;
        RECT 10.750 0.580 11.680 0.750 ;
        RECT 10.750 0.535 10.920 0.580 ;
        RECT 9.385 0.365 10.920 0.535 ;
        RECT 11.935 0.425 12.265 0.960 ;
        RECT 12.465 0.790 13.565 0.960 ;
        RECT 12.465 0.595 12.795 0.790 ;
        RECT 12.975 0.425 13.225 0.620 ;
        RECT 11.415 0.085 11.755 0.410 ;
        RECT 11.935 0.255 13.225 0.425 ;
        RECT 13.395 0.500 13.565 0.790 ;
        RECT 13.735 0.670 13.905 1.130 ;
        RECT 14.550 1.020 14.720 1.300 ;
        RECT 14.075 0.850 14.720 1.020 ;
        RECT 15.450 1.220 16.375 1.550 ;
        RECT 14.075 0.500 14.245 0.850 ;
        RECT 13.395 0.330 14.245 0.500 ;
        RECT 14.415 0.085 14.735 0.680 ;
        RECT 15.450 0.350 15.725 1.220 ;
        RECT 15.905 0.085 16.155 1.050 ;
        RECT 0.000 -0.085 16.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 5.435 1.580 5.605 1.750 ;
        RECT 8.315 1.950 8.485 2.120 ;
        RECT 9.755 1.580 9.925 1.750 ;
        RECT 11.675 1.950 11.845 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
      LAYER met1 ;
        RECT 5.375 1.735 5.665 1.780 ;
        RECT 9.695 1.735 9.985 1.780 ;
        RECT 5.375 1.595 9.985 1.735 ;
        RECT 5.375 1.550 5.665 1.595 ;
        RECT 9.695 1.550 9.985 1.595 ;
  END
END sky130_fd_sc_hs__sdfbbn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfbbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.240 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.350 3.895 1.780 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.460 1.815 1.790 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 13.945 1.505 14.275 1.835 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.125 0.550 2.135 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.125 1.315 1.795 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER met1 ;
        RECT 9.215 1.735 9.505 1.780 ;
        RECT 12.095 1.735 12.385 1.780 ;
        RECT 9.215 1.595 12.385 1.735 ;
        RECT 9.215 1.550 9.505 1.595 ;
        RECT 12.095 1.550 12.385 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 18.240 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.310 1.175 5.130 1.360 ;
        RECT 7.235 1.175 9.890 1.305 ;
        RECT 13.715 1.240 14.655 1.450 ;
        RECT 3.310 1.145 9.890 1.175 ;
        RECT 0.030 1.090 9.890 1.145 ;
        RECT 0.030 0.960 10.365 1.090 ;
        RECT 11.730 0.960 18.235 1.240 ;
        RECT 0.030 0.245 18.235 0.960 ;
        RECT 0.000 0.000 18.240 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 18.430 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 18.240 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 17.395 1.820 17.705 2.980 ;
        RECT 17.535 1.050 17.705 1.820 ;
        RECT 17.370 0.350 17.705 1.050 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 15.375 1.780 15.625 2.980 ;
        RECT 15.375 1.550 15.715 1.780 ;
        RECT 15.375 1.220 15.610 1.550 ;
        RECT 15.280 0.350 15.610 1.220 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 18.240 3.415 ;
        RECT 0.115 2.475 0.365 2.980 ;
        RECT 0.565 2.645 0.895 3.245 ;
        RECT 1.065 2.905 2.185 3.075 ;
        RECT 1.065 2.475 1.235 2.905 ;
        RECT 0.115 2.305 1.235 2.475 ;
        RECT 1.405 2.300 1.655 2.735 ;
        RECT 1.855 2.300 2.185 2.905 ;
        RECT 2.415 2.300 2.745 3.245 ;
        RECT 1.485 2.130 1.655 2.300 ;
        RECT 1.485 1.960 2.155 2.130 ;
        RECT 1.985 1.290 2.155 1.960 ;
        RECT 2.945 1.810 3.195 2.980 ;
        RECT 3.425 2.120 3.675 2.980 ;
        RECT 3.875 2.290 4.205 3.245 ;
        RECT 3.425 1.950 4.235 2.120 ;
        RECT 2.605 1.480 3.195 1.810 ;
        RECT 1.485 1.120 2.770 1.290 ;
        RECT 1.485 0.955 1.690 1.120 ;
        RECT 0.140 0.085 0.470 0.955 ;
        RECT 0.960 0.625 1.690 0.955 ;
        RECT 2.180 0.085 2.430 0.950 ;
        RECT 2.600 0.425 2.770 1.120 ;
        RECT 2.940 0.595 3.195 1.480 ;
        RECT 4.065 1.670 4.235 1.950 ;
        RECT 4.405 1.840 4.785 2.980 ;
        RECT 4.965 2.350 5.215 3.245 ;
        RECT 5.385 2.905 7.825 3.075 ;
        RECT 5.385 2.180 5.555 2.905 ;
        RECT 6.900 2.900 7.825 2.905 ;
        RECT 4.065 1.340 4.445 1.670 ;
        RECT 4.615 1.350 4.785 1.840 ;
        RECT 5.035 2.010 5.555 2.180 ;
        RECT 5.840 2.210 6.170 2.735 ;
        RECT 6.340 2.550 6.670 2.735 ;
        RECT 6.900 2.730 8.045 2.900 ;
        RECT 6.340 2.380 7.705 2.550 ;
        RECT 5.840 2.040 7.365 2.210 ;
        RECT 5.035 1.830 5.365 2.010 ;
        RECT 6.495 1.840 6.825 1.855 ;
        RECT 5.595 1.525 6.825 1.840 ;
        RECT 5.595 1.350 6.115 1.525 ;
        RECT 7.035 1.355 7.365 2.040 ;
        RECT 4.065 1.170 4.235 1.340 ;
        RECT 4.615 1.180 6.115 1.350 ;
        RECT 6.285 1.185 7.365 1.355 ;
        RECT 3.420 1.000 4.235 1.170 ;
        RECT 3.365 0.660 4.520 0.830 ;
        RECT 3.365 0.425 3.535 0.660 ;
        RECT 2.600 0.255 3.535 0.425 ;
        RECT 3.930 0.085 4.180 0.490 ;
        RECT 4.350 0.425 4.520 0.660 ;
        RECT 4.690 0.595 4.940 1.180 ;
        RECT 5.110 0.840 6.115 1.010 ;
        RECT 5.110 0.425 5.280 0.840 ;
        RECT 4.350 0.255 5.280 0.425 ;
        RECT 5.450 0.085 5.720 0.670 ;
        RECT 5.945 0.435 6.115 0.840 ;
        RECT 6.285 0.605 6.615 1.185 ;
        RECT 7.535 1.015 7.705 2.380 ;
        RECT 6.785 0.845 7.705 1.015 ;
        RECT 7.875 2.295 8.045 2.730 ;
        RECT 8.365 2.465 8.695 3.245 ;
        RECT 8.905 2.295 9.235 2.980 ;
        RECT 7.875 2.125 9.235 2.295 ;
        RECT 9.465 2.290 9.795 3.245 ;
        RECT 7.875 1.115 8.045 2.125 ;
        RECT 8.905 2.120 9.235 2.125 ;
        RECT 10.305 2.270 10.635 2.980 ;
        RECT 11.230 2.600 11.560 3.245 ;
        RECT 11.805 2.430 12.135 2.980 ;
        RECT 12.305 2.600 12.635 3.245 ;
        RECT 13.185 2.675 13.435 2.980 ;
        RECT 14.280 2.845 15.170 3.245 ;
        RECT 13.185 2.505 14.655 2.675 ;
        RECT 13.185 2.430 13.435 2.505 ;
        RECT 8.215 1.285 8.620 1.955 ;
        RECT 8.905 1.950 9.945 2.120 ;
        RECT 10.305 2.100 10.910 2.270 ;
        RECT 8.790 1.450 9.445 1.780 ;
        RECT 9.615 1.580 9.945 1.950 ;
        RECT 10.740 1.920 10.910 2.100 ;
        RECT 11.080 2.260 13.435 2.430 ;
        RECT 11.080 2.090 11.410 2.260 ;
        RECT 11.580 1.920 12.665 2.090 ;
        RECT 13.185 2.060 13.435 2.260 ;
        RECT 10.155 1.580 10.485 1.755 ;
        RECT 10.740 1.750 11.750 1.920 ;
        RECT 12.495 1.890 12.665 1.920 ;
        RECT 13.605 2.005 14.075 2.335 ;
        RECT 8.450 1.280 8.620 1.285 ;
        RECT 10.155 1.280 11.385 1.580 ;
        RECT 7.875 0.945 8.280 1.115 ;
        RECT 8.450 1.110 9.725 1.280 ;
        RECT 10.155 1.180 10.485 1.280 ;
        RECT 11.555 1.110 11.725 1.750 ;
        RECT 11.955 1.180 12.325 1.750 ;
        RECT 12.495 1.720 13.365 1.890 ;
        RECT 12.495 1.300 12.825 1.550 ;
        RECT 13.035 1.470 13.365 1.720 ;
        RECT 13.605 1.335 13.775 2.005 ;
        RECT 14.485 1.760 14.655 2.505 ;
        RECT 14.825 1.950 15.170 2.845 ;
        RECT 15.825 1.950 16.155 3.245 ;
        RECT 14.485 1.430 14.815 1.760 ;
        RECT 16.340 1.550 16.700 2.940 ;
        RECT 16.895 1.820 17.225 3.245 ;
        RECT 17.875 1.820 18.125 3.245 ;
        RECT 13.605 1.300 14.150 1.335 ;
        RECT 6.785 0.435 7.115 0.845 ;
        RECT 5.945 0.265 7.115 0.435 ;
        RECT 7.345 0.435 7.770 0.675 ;
        RECT 7.950 0.605 8.280 0.945 ;
        RECT 8.450 0.605 8.885 0.935 ;
        RECT 8.450 0.435 8.620 0.605 ;
        RECT 7.345 0.265 8.620 0.435 ;
        RECT 9.055 0.085 9.385 0.940 ;
        RECT 9.555 0.430 9.725 1.110 ;
        RECT 10.940 0.940 11.725 1.110 ;
        RECT 12.495 1.130 14.150 1.300 ;
        RECT 12.495 0.940 12.665 1.130 ;
        RECT 13.605 1.005 14.150 1.130 ;
        RECT 14.485 1.005 14.655 1.430 ;
        RECT 16.340 1.220 17.365 1.550 ;
        RECT 10.940 0.850 11.110 0.940 ;
        RECT 9.960 0.600 11.110 0.850 ;
        RECT 11.895 0.770 12.665 0.940 ;
        RECT 12.835 0.835 13.085 0.960 ;
        RECT 14.320 0.835 14.655 1.005 ;
        RECT 11.340 0.600 12.065 0.770 ;
        RECT 12.835 0.665 14.490 0.835 ;
        RECT 11.340 0.430 11.510 0.600 ;
        RECT 9.555 0.260 11.510 0.430 ;
        RECT 11.680 0.085 12.055 0.430 ;
        RECT 12.235 0.425 12.655 0.600 ;
        RECT 12.835 0.595 13.085 0.665 ;
        RECT 13.265 0.425 13.595 0.495 ;
        RECT 12.235 0.255 13.595 0.425 ;
        RECT 14.825 0.085 15.110 1.130 ;
        RECT 15.780 0.085 16.110 1.130 ;
        RECT 16.340 0.540 16.670 1.220 ;
        RECT 16.870 0.085 17.200 1.050 ;
        RECT 17.880 0.085 18.130 1.130 ;
        RECT 0.000 -0.085 18.240 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 16.955 3.245 17.125 3.415 ;
        RECT 17.435 3.245 17.605 3.415 ;
        RECT 17.915 3.245 18.085 3.415 ;
        RECT 5.915 1.210 6.085 1.380 ;
        RECT 9.275 1.580 9.445 1.750 ;
        RECT 10.235 1.210 10.405 1.380 ;
        RECT 12.155 1.580 12.325 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
        RECT 17.435 -0.085 17.605 0.085 ;
        RECT 17.915 -0.085 18.085 0.085 ;
      LAYER met1 ;
        RECT 5.855 1.365 6.145 1.410 ;
        RECT 10.175 1.365 10.465 1.410 ;
        RECT 5.855 1.225 10.465 1.365 ;
        RECT 5.855 1.180 6.145 1.225 ;
        RECT 10.175 1.180 10.465 1.225 ;
  END
END sky130_fd_sc_hs__sdfbbn_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfbbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.430 1.180 3.760 1.670 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.525 1.765 1.855 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 13.065 1.180 13.360 1.550 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.125 0.550 2.135 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.550 1.285 2.095 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER li1 ;
        RECT 7.095 2.905 8.105 3.075 ;
        RECT 7.095 1.655 7.265 2.905 ;
        RECT 7.935 2.335 8.105 2.905 ;
        RECT 8.855 2.905 10.265 3.075 ;
        RECT 8.855 2.335 9.025 2.905 ;
        RECT 7.935 2.165 9.025 2.335 ;
        RECT 10.095 2.185 10.265 2.905 ;
        RECT 10.095 2.015 10.295 2.185 ;
        RECT 10.125 1.860 10.295 2.015 ;
        RECT 11.055 1.860 11.365 2.150 ;
        RECT 10.125 1.800 11.365 1.860 ;
        RECT 10.125 1.690 11.385 1.800 ;
        RECT 7.045 1.410 7.375 1.655 ;
        RECT 11.055 1.520 11.385 1.690 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 15.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.980 1.145 4.855 1.360 ;
        RECT 6.560 1.275 7.470 1.305 ;
        RECT 6.560 1.240 10.175 1.275 ;
        RECT 6.560 1.175 15.835 1.240 ;
        RECT 0.030 1.030 4.855 1.145 ;
        RECT 5.905 1.030 15.835 1.175 ;
        RECT 0.030 0.245 15.835 1.030 ;
        RECT 0.000 0.000 15.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.030 3.520 ;
        RECT 12.680 1.560 14.260 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 15.840 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 15.395 0.350 15.735 2.980 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518900 ;
    PORT
      LAYER li1 ;
        RECT 13.870 1.720 14.275 2.890 ;
        RECT 14.105 1.050 14.275 1.720 ;
        RECT 13.770 0.350 14.275 1.050 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 15.840 3.415 ;
        RECT 0.115 2.475 0.445 2.980 ;
        RECT 0.615 2.645 0.945 3.245 ;
        RECT 1.115 2.905 2.275 3.075 ;
        RECT 1.115 2.475 1.285 2.905 ;
        RECT 0.115 2.305 1.285 2.475 ;
        RECT 1.495 2.195 1.745 2.735 ;
        RECT 1.945 2.520 2.275 2.905 ;
        RECT 2.505 2.520 2.755 3.245 ;
        RECT 2.955 2.350 3.285 2.980 ;
        RECT 1.495 2.025 2.105 2.195 ;
        RECT 1.935 1.355 2.105 2.025 ;
        RECT 2.275 2.180 3.285 2.350 ;
        RECT 2.275 1.830 2.780 2.180 ;
        RECT 3.515 2.010 3.845 2.980 ;
        RECT 4.045 2.180 4.215 3.245 ;
        RECT 1.040 1.185 2.420 1.355 ;
        RECT 0.140 0.085 0.470 0.955 ;
        RECT 1.040 0.575 1.370 1.185 ;
        RECT 1.830 0.085 2.080 1.015 ;
        RECT 2.250 0.425 2.420 1.185 ;
        RECT 2.610 1.035 2.780 1.830 ;
        RECT 3.090 1.840 4.245 2.010 ;
        RECT 4.415 1.840 4.905 2.980 ;
        RECT 5.075 2.035 5.405 2.755 ;
        RECT 5.575 2.205 6.125 2.535 ;
        RECT 5.075 1.865 5.785 2.035 ;
        RECT 2.610 0.595 2.860 1.035 ;
        RECT 3.090 1.010 3.260 1.840 ;
        RECT 4.075 1.670 4.245 1.840 ;
        RECT 4.735 1.695 4.905 1.840 ;
        RECT 4.075 1.340 4.565 1.670 ;
        RECT 4.735 1.365 5.445 1.695 ;
        RECT 4.735 1.170 4.905 1.365 ;
        RECT 5.615 1.195 5.785 1.865 ;
        RECT 3.090 0.595 3.340 1.010 ;
        RECT 4.360 1.000 4.905 1.170 ;
        RECT 5.165 1.025 5.785 1.195 ;
        RECT 5.955 1.825 6.125 2.205 ;
        RECT 6.595 2.075 6.925 3.245 ;
        RECT 7.435 1.995 7.765 2.735 ;
        RECT 8.315 2.505 8.685 3.245 ;
        RECT 9.375 2.110 9.925 2.735 ;
        RECT 10.435 2.660 11.150 3.245 ;
        RECT 11.535 2.490 11.785 2.980 ;
        RECT 7.435 1.825 9.015 1.995 ;
        RECT 5.955 1.655 6.875 1.825 ;
        RECT 5.165 0.830 5.335 1.025 ;
        RECT 5.955 0.855 6.125 1.655 ;
        RECT 3.510 0.660 5.335 0.830 ;
        RECT 3.510 0.425 3.680 0.660 ;
        RECT 2.250 0.255 3.680 0.425 ;
        RECT 3.850 0.085 4.180 0.490 ;
        RECT 5.005 0.460 5.335 0.660 ;
        RECT 5.505 0.685 6.125 0.855 ;
        RECT 6.295 0.900 6.535 1.485 ;
        RECT 6.705 1.240 6.875 1.655 ;
        RECT 7.585 1.240 7.915 1.585 ;
        RECT 6.705 1.070 7.915 1.240 ;
        RECT 8.125 1.180 8.515 1.585 ;
        RECT 8.685 1.335 9.015 1.825 ;
        RECT 9.255 1.505 9.585 1.940 ;
        RECT 9.755 1.845 9.925 2.110 ;
        RECT 10.465 2.320 11.785 2.490 ;
        RECT 12.295 2.480 12.625 3.245 ;
        RECT 13.340 2.480 13.670 3.245 ;
        RECT 10.465 2.030 10.795 2.320 ;
        RECT 11.535 2.310 11.785 2.320 ;
        RECT 11.535 2.140 13.700 2.310 ;
        RECT 11.535 1.970 12.215 2.140 ;
        RECT 9.755 1.675 9.955 1.845 ;
        RECT 9.785 1.520 9.955 1.675 ;
        RECT 9.255 1.335 9.615 1.505 ;
        RECT 8.685 0.900 8.855 1.335 ;
        RECT 6.295 0.730 8.855 0.900 ;
        RECT 5.505 0.460 5.835 0.685 ;
        RECT 7.820 0.655 8.150 0.730 ;
        RECT 6.490 0.085 6.885 0.560 ;
        RECT 7.145 0.480 7.640 0.560 ;
        RECT 8.330 0.480 8.715 0.560 ;
        RECT 7.145 0.310 8.715 0.480 ;
        RECT 9.025 0.085 9.275 1.050 ;
        RECT 9.445 0.425 9.615 1.335 ;
        RECT 9.785 1.350 10.885 1.520 ;
        RECT 11.595 1.350 11.875 1.550 ;
        RECT 9.785 0.595 9.985 1.350 ;
        RECT 10.715 1.180 11.875 1.350 ;
        RECT 10.155 0.425 10.485 1.180 ;
        RECT 12.045 1.010 12.215 1.970 ;
        RECT 12.725 1.720 13.155 1.970 ;
        RECT 12.445 1.180 12.895 1.720 ;
        RECT 13.530 1.550 13.700 2.140 ;
        RECT 14.445 1.685 14.775 2.980 ;
        RECT 14.945 2.115 15.205 3.245 ;
        RECT 13.530 1.220 13.915 1.550 ;
        RECT 14.445 1.355 14.845 1.685 ;
        RECT 12.725 1.010 12.895 1.180 ;
        RECT 9.445 0.255 10.485 0.425 ;
        RECT 10.900 0.085 11.150 1.010 ;
        RECT 11.330 0.425 11.660 1.010 ;
        RECT 11.870 0.595 12.215 1.010 ;
        RECT 12.385 0.425 12.555 1.010 ;
        RECT 12.725 0.670 13.115 1.010 ;
        RECT 11.330 0.255 12.555 0.425 ;
        RECT 13.295 0.085 13.590 1.000 ;
        RECT 14.445 0.350 14.715 1.355 ;
        RECT 14.895 0.085 15.225 0.940 ;
        RECT 0.000 -0.085 15.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 8.315 1.210 8.485 1.380 ;
        RECT 12.635 1.210 12.805 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
      LAYER met1 ;
        RECT 8.255 1.365 8.545 1.410 ;
        RECT 12.575 1.365 12.865 1.410 ;
        RECT 8.255 1.225 12.865 1.365 ;
        RECT 8.255 1.180 8.545 1.225 ;
        RECT 12.575 1.180 12.865 1.225 ;
  END
END sky130_fd_sc_hs__sdfbbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.180 4.645 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.810 2.100 1.310 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 3.935 2.105 4.225 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 10.655 2.105 10.945 2.150 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 3.935 1.920 4.225 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
        RECT 10.655 1.920 10.945 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.935 1.440 3.265 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.660 1.795 1.880 ;
        RECT 0.605 1.490 2.725 1.660 ;
        RECT 2.395 1.260 2.725 1.490 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.120 1.035 5.530 1.240 ;
        RECT 7.775 1.035 9.115 1.140 ;
        RECT 2.160 1.000 9.115 1.035 ;
        RECT 0.995 0.920 9.115 1.000 ;
        RECT 11.405 0.920 13.910 1.240 ;
        RECT 0.005 0.245 13.910 0.920 ;
        RECT 0.000 0.000 13.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.110 3.520 ;
        RECT 4.095 1.640 9.515 1.660 ;
        RECT 8.005 1.555 9.515 1.640 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.920 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518900 ;
    PORT
      LAYER li1 ;
        RECT 13.555 1.820 13.835 2.980 ;
        RECT 13.665 1.130 13.835 1.820 ;
        RECT 13.470 0.350 13.835 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.537600 ;
    PORT
      LAYER li1 ;
        RECT 12.015 0.350 12.345 2.980 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.920 3.415 ;
        RECT 0.115 2.220 1.055 2.975 ;
        RECT 1.225 2.390 1.555 3.245 ;
        RECT 2.095 2.560 2.425 3.000 ;
        RECT 3.085 2.730 3.445 3.245 ;
        RECT 3.615 2.560 3.985 3.000 ;
        RECT 4.705 2.690 5.035 3.245 ;
        RECT 2.095 2.520 3.985 2.560 ;
        RECT 5.725 2.520 5.975 2.755 ;
        RECT 2.095 2.390 5.975 2.520 ;
        RECT 6.175 2.490 6.845 2.755 ;
        RECT 7.090 2.660 7.420 3.245 ;
        RECT 7.615 2.490 7.945 2.755 ;
        RECT 6.175 2.415 7.945 2.490 ;
        RECT 3.445 2.350 5.975 2.390 ;
        RECT 3.445 2.320 3.985 2.350 ;
        RECT 0.115 2.050 2.695 2.220 ;
        RECT 0.115 1.310 0.285 2.050 ;
        RECT 2.365 1.830 2.695 2.050 ;
        RECT 0.115 0.980 1.395 1.310 ;
        RECT 3.445 1.090 3.615 2.320 ;
        RECT 5.725 2.300 5.975 2.350 ;
        RECT 5.805 2.245 5.975 2.300 ;
        RECT 6.675 2.320 7.945 2.415 ;
        RECT 3.785 1.820 4.165 2.150 ;
        RECT 4.335 1.970 4.585 2.180 ;
        RECT 4.335 1.800 4.985 1.970 ;
        RECT 5.155 1.905 5.620 2.130 ;
        RECT 5.805 2.075 6.505 2.245 ;
        RECT 5.155 1.800 6.165 1.905 ;
        RECT 0.115 0.350 0.365 0.980 ;
        RECT 2.270 0.920 3.615 1.090 ;
        RECT 4.815 1.630 4.985 1.800 ;
        RECT 4.815 1.300 5.280 1.630 ;
        RECT 5.450 1.575 6.165 1.800 ;
        RECT 4.815 1.010 4.985 1.300 ;
        RECT 5.450 1.130 5.620 1.575 ;
        RECT 6.335 1.265 6.505 2.075 ;
        RECT 0.545 0.085 0.875 0.810 ;
        RECT 1.105 0.425 1.355 0.810 ;
        RECT 2.270 0.595 2.600 0.920 ;
        RECT 4.230 0.840 4.985 1.010 ;
        RECT 5.170 0.960 5.620 1.130 ;
        RECT 5.810 1.095 6.505 1.265 ;
        RECT 3.170 0.425 3.500 0.750 ;
        RECT 1.105 0.255 3.500 0.425 ;
        RECT 3.670 0.085 4.000 0.750 ;
        RECT 4.230 0.350 4.480 0.840 ;
        RECT 4.660 0.085 4.990 0.670 ;
        RECT 5.170 0.425 5.420 0.960 ;
        RECT 5.810 0.790 5.980 1.095 ;
        RECT 6.675 0.925 6.845 2.320 ;
        RECT 7.015 1.105 7.235 1.760 ;
        RECT 7.405 1.545 7.575 2.320 ;
        RECT 7.745 1.820 8.035 2.150 ;
        RECT 8.235 1.715 8.485 3.245 ;
        RECT 7.405 1.275 8.270 1.545 ;
        RECT 8.685 1.415 8.935 2.755 ;
        RECT 9.105 2.425 10.095 2.755 ;
        RECT 10.305 2.660 10.650 3.245 ;
        RECT 10.855 2.490 11.185 2.885 ;
        RECT 11.370 2.695 11.815 3.245 ;
        RECT 9.105 1.755 9.325 2.425 ;
        RECT 9.505 1.575 9.755 2.230 ;
        RECT 8.440 1.245 8.935 1.415 ;
        RECT 9.105 1.345 9.755 1.575 ;
        RECT 9.925 1.435 10.095 2.425 ;
        RECT 10.265 2.320 11.405 2.490 ;
        RECT 10.265 1.650 10.525 2.320 ;
        RECT 10.695 1.685 11.065 2.150 ;
        RECT 11.235 1.800 11.405 2.320 ;
        RECT 11.585 1.970 11.815 2.695 ;
        RECT 11.235 1.630 11.845 1.800 ;
        RECT 8.440 1.105 8.610 1.245 ;
        RECT 7.015 0.935 8.610 1.105 ;
        RECT 9.105 1.075 9.435 1.345 ;
        RECT 9.925 1.175 11.425 1.435 ;
        RECT 5.650 0.595 5.980 0.790 ;
        RECT 6.150 0.595 6.845 0.925 ;
        RECT 7.015 0.595 8.110 0.765 ;
        RECT 8.280 0.595 8.610 0.935 ;
        RECT 8.780 0.905 9.435 1.075 ;
        RECT 9.605 1.005 11.425 1.175 ;
        RECT 7.015 0.425 7.185 0.595 ;
        RECT 7.940 0.425 8.110 0.595 ;
        RECT 8.780 0.425 8.950 0.905 ;
        RECT 9.605 0.735 9.775 1.005 ;
        RECT 5.170 0.255 7.185 0.425 ;
        RECT 7.440 0.085 7.770 0.425 ;
        RECT 7.940 0.255 8.950 0.425 ;
        RECT 9.135 0.405 9.775 0.735 ;
        RECT 10.165 0.085 10.495 0.760 ;
        RECT 11.675 0.750 11.845 1.630 ;
        RECT 10.955 0.580 11.845 0.750 ;
        RECT 12.570 1.630 12.855 2.980 ;
        RECT 13.045 1.820 13.325 3.245 ;
        RECT 12.570 1.300 13.485 1.630 ;
        RECT 10.955 0.350 11.285 0.580 ;
        RECT 12.570 0.455 12.855 1.300 ;
        RECT 11.510 0.085 11.840 0.410 ;
        RECT 13.120 0.085 13.290 1.130 ;
        RECT 0.000 -0.085 13.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 10.715 1.950 10.885 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
  END
END sky130_fd_sc_hs__sdfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.880 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.905 1.180 4.235 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.810 2.090 1.190 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 3.935 2.105 4.225 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 10.655 2.105 10.945 2.150 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 3.935 1.920 4.225 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
        RECT 10.655 1.920 10.945 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.440 3.275 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.540 1.820 1.795 2.150 ;
        RECT 1.625 1.620 1.795 1.820 ;
        RECT 1.625 1.360 2.735 1.620 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.130 1.140 5.540 1.240 ;
        RECT 4.130 0.945 9.330 1.140 ;
        RECT 0.005 0.920 9.330 0.945 ;
        RECT 11.555 0.920 14.875 1.240 ;
        RECT 0.005 0.245 14.875 0.920 ;
        RECT 0.000 0.000 14.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 15.070 3.520 ;
        RECT 7.970 1.595 12.540 1.660 ;
        RECT 7.970 1.555 9.470 1.595 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.880 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 14.055 0.350 14.325 2.980 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 12.030 1.085 12.360 2.980 ;
        RECT 12.030 0.915 12.465 1.085 ;
        RECT 12.135 0.350 12.465 0.915 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.880 3.415 ;
        RECT 0.115 2.490 0.445 2.980 ;
        RECT 0.615 2.730 1.400 3.245 ;
        RECT 1.940 2.660 2.945 2.910 ;
        RECT 3.115 2.660 3.445 3.245 ;
        RECT 2.775 2.490 2.945 2.660 ;
        RECT 3.615 2.520 3.995 2.980 ;
        RECT 4.705 2.690 5.035 3.245 ;
        RECT 5.710 2.520 5.985 2.725 ;
        RECT 3.615 2.490 5.985 2.520 ;
        RECT 0.115 2.320 2.605 2.490 ;
        RECT 2.775 2.350 5.985 2.490 ;
        RECT 2.775 2.320 3.995 2.350 ;
        RECT 5.710 2.330 5.985 2.350 ;
        RECT 6.160 2.510 6.660 2.725 ;
        RECT 7.070 2.680 7.320 3.245 ;
        RECT 7.550 2.510 7.915 2.725 ;
        RECT 6.160 2.340 7.915 2.510 ;
        RECT 0.115 1.580 0.285 2.320 ;
        RECT 2.275 1.830 2.605 2.320 ;
        RECT 0.115 1.250 1.395 1.580 ;
        RECT 0.115 0.375 0.365 1.250 ;
        RECT 3.445 1.175 3.615 2.320 ;
        RECT 3.785 1.820 4.165 2.150 ;
        RECT 4.335 1.990 4.585 2.180 ;
        RECT 5.815 2.170 5.985 2.330 ;
        RECT 4.335 1.820 4.985 1.990 ;
        RECT 5.155 1.830 5.645 2.160 ;
        RECT 5.815 2.000 6.490 2.170 ;
        RECT 4.815 1.660 4.985 1.820 ;
        RECT 4.815 1.500 5.305 1.660 ;
        RECT 2.260 1.005 3.615 1.175 ;
        RECT 4.405 1.330 5.305 1.500 ;
        RECT 5.475 1.500 6.150 1.830 ;
        RECT 4.405 1.010 4.575 1.330 ;
        RECT 5.475 1.160 5.645 1.500 ;
        RECT 6.320 1.290 6.490 2.000 ;
        RECT 0.545 0.085 0.875 0.835 ;
        RECT 1.095 0.425 1.345 0.835 ;
        RECT 2.260 0.595 2.610 1.005 ;
        RECT 3.100 0.425 3.430 0.835 ;
        RECT 1.095 0.255 3.430 0.425 ;
        RECT 3.640 0.085 3.970 0.835 ;
        RECT 4.240 0.350 4.575 1.010 ;
        RECT 4.750 0.085 4.920 1.130 ;
        RECT 5.100 0.990 5.645 1.160 ;
        RECT 5.820 1.120 6.490 1.290 ;
        RECT 5.100 0.480 5.430 0.990 ;
        RECT 5.820 0.820 5.990 1.120 ;
        RECT 6.660 0.950 6.830 2.340 ;
        RECT 7.380 2.320 7.915 2.340 ;
        RECT 5.660 0.650 5.990 0.820 ;
        RECT 6.160 0.650 6.830 0.950 ;
        RECT 7.000 1.090 7.210 1.775 ;
        RECT 7.380 1.575 7.550 2.320 ;
        RECT 7.720 1.795 8.020 2.150 ;
        RECT 8.190 1.745 8.440 3.245 ;
        RECT 8.640 1.745 8.930 2.755 ;
        RECT 9.100 2.365 10.095 2.695 ;
        RECT 10.265 2.660 10.860 3.245 ;
        RECT 11.065 2.490 11.395 2.795 ;
        RECT 7.380 1.260 8.590 1.575 ;
        RECT 8.760 1.090 8.930 1.745 ;
        RECT 9.310 1.865 9.755 2.195 ;
        RECT 9.310 1.235 9.640 1.865 ;
        RECT 7.000 0.920 8.930 1.090 ;
        RECT 7.000 0.580 8.325 0.750 ;
        RECT 8.495 0.595 8.930 0.920 ;
        RECT 9.100 0.905 9.640 1.235 ;
        RECT 9.925 1.310 10.095 2.365 ;
        RECT 10.265 2.320 11.395 2.490 ;
        RECT 10.265 1.650 10.545 2.320 ;
        RECT 10.715 1.820 11.395 2.150 ;
        RECT 11.600 1.820 11.850 3.245 ;
        RECT 12.540 1.920 12.830 3.245 ;
        RECT 10.265 1.480 11.860 1.650 ;
        RECT 9.925 1.045 11.520 1.310 ;
        RECT 7.000 0.480 7.170 0.580 ;
        RECT 5.100 0.310 7.170 0.480 ;
        RECT 8.155 0.425 8.325 0.580 ;
        RECT 9.100 0.425 9.270 0.905 ;
        RECT 9.925 0.735 10.095 1.045 ;
        RECT 11.690 0.875 11.860 1.480 ;
        RECT 13.065 1.630 13.325 2.980 ;
        RECT 13.545 1.820 13.875 3.245 ;
        RECT 14.495 1.820 14.775 3.245 ;
        RECT 13.065 1.300 13.885 1.630 ;
        RECT 7.450 0.085 7.985 0.410 ;
        RECT 8.155 0.255 9.270 0.425 ;
        RECT 9.440 0.405 10.095 0.735 ;
        RECT 10.335 0.085 10.665 0.810 ;
        RECT 11.125 0.705 11.860 0.875 ;
        RECT 11.125 0.350 11.455 0.705 ;
        RECT 11.645 0.085 11.895 0.535 ;
        RECT 12.635 0.085 12.895 1.050 ;
        RECT 13.065 0.350 13.325 1.300 ;
        RECT 13.670 0.085 13.840 1.130 ;
        RECT 14.495 0.085 14.780 1.130 ;
        RECT 0.000 -0.085 14.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 10.715 1.950 10.885 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
  END
END sky130_fd_sc_hs__sdfrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.210 4.675 1.550 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.780 1.980 2.120 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 3.455 1.735 3.745 1.780 ;
        RECT 7.775 1.735 8.065 1.780 ;
        RECT 11.135 1.735 11.425 1.780 ;
        RECT 3.455 1.595 11.425 1.735 ;
        RECT 3.455 1.550 3.745 1.595 ;
        RECT 7.775 1.550 8.065 1.595 ;
        RECT 11.135 1.550 11.425 1.595 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.800 1.525 3.235 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.580 0.865 2.080 ;
        RECT 0.535 1.410 2.045 1.580 ;
        RECT 1.875 0.955 2.550 1.410 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.695 1.240 5.785 1.310 ;
        RECT 3.740 1.205 5.785 1.240 ;
        RECT 7.895 1.205 9.515 1.490 ;
        RECT 0.005 0.955 1.055 0.990 ;
        RECT 3.740 0.955 9.515 1.205 ;
        RECT 12.865 1.050 13.915 1.240 ;
        RECT 0.005 0.920 9.515 0.955 ;
        RECT 12.355 0.920 13.915 1.050 ;
        RECT 0.005 0.245 13.915 0.920 ;
        RECT 0.000 0.000 13.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.780 14.110 3.520 ;
        RECT -0.190 1.660 5.995 1.780 ;
        RECT 9.725 1.660 14.110 1.780 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.920 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.546900 ;
    PORT
      LAYER li1 ;
        RECT 13.475 0.350 13.805 2.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.920 3.415 ;
        RECT 0.115 2.460 0.365 2.980 ;
        RECT 0.565 2.630 0.895 3.245 ;
        RECT 2.815 2.970 3.145 3.245 ;
        RECT 1.405 2.800 2.220 2.960 ;
        RECT 3.430 2.800 3.680 2.980 ;
        RECT 1.405 2.630 3.680 2.800 ;
        RECT 3.910 2.645 4.240 3.245 ;
        RECT 4.995 2.645 5.325 3.245 ;
        RECT 3.430 2.475 3.680 2.630 ;
        RECT 6.005 2.475 6.255 2.980 ;
        RECT 0.115 2.290 2.545 2.460 ;
        RECT 3.430 2.305 6.255 2.475 ;
        RECT 6.455 2.445 6.785 2.980 ;
        RECT 7.295 2.615 7.545 3.245 ;
        RECT 7.745 2.445 8.075 2.980 ;
        RECT 3.430 2.300 4.075 2.305 ;
        RECT 0.115 1.240 0.365 2.290 ;
        RECT 2.215 1.580 2.545 2.290 ;
        RECT 3.405 1.355 3.735 2.025 ;
        RECT 0.115 1.050 1.620 1.240 ;
        RECT 3.905 1.185 4.075 2.300 ;
        RECT 6.455 2.275 8.075 2.445 ;
        RECT 8.295 2.310 8.625 3.245 ;
        RECT 4.435 1.820 5.015 2.135 ;
        RECT 0.115 0.420 0.445 1.050 ;
        RECT 1.290 0.935 1.620 1.050 ;
        RECT 2.720 1.015 4.075 1.185 ;
        RECT 4.845 1.620 5.015 1.820 ;
        RECT 5.345 2.105 5.775 2.135 ;
        RECT 5.345 1.820 6.590 2.105 ;
        RECT 4.845 1.290 5.175 1.620 ;
        RECT 5.345 1.435 5.675 1.820 ;
        RECT 6.260 1.775 6.590 1.820 ;
        RECT 4.845 1.040 5.015 1.290 ;
        RECT 0.615 0.085 0.945 0.880 ;
        RECT 2.720 0.765 2.890 1.015 ;
        RECT 1.165 0.425 1.495 0.765 ;
        RECT 1.955 0.595 2.890 0.765 ;
        RECT 3.060 0.425 3.390 0.845 ;
        RECT 3.905 0.700 4.075 1.015 ;
        RECT 4.245 0.870 5.015 1.040 ;
        RECT 5.345 1.265 6.495 1.435 ;
        RECT 5.345 0.870 5.675 1.265 ;
        RECT 5.905 0.700 6.155 1.095 ;
        RECT 3.905 0.530 6.155 0.700 ;
        RECT 6.325 0.545 6.495 1.265 ;
        RECT 6.760 1.095 6.930 2.275 ;
        RECT 7.905 2.140 8.075 2.275 ;
        RECT 8.795 2.140 9.565 2.980 ;
        RECT 7.905 1.970 8.520 2.140 ;
        RECT 7.145 1.300 7.475 1.870 ;
        RECT 7.685 1.470 8.035 1.800 ;
        RECT 8.225 1.470 8.520 1.970 ;
        RECT 8.690 1.970 9.565 2.140 ;
        RECT 8.690 1.300 8.860 1.970 ;
        RECT 9.735 1.880 10.065 2.980 ;
        RECT 10.605 2.650 11.210 3.245 ;
        RECT 11.380 2.460 11.710 2.980 ;
        RECT 11.880 2.630 12.210 3.245 ;
        RECT 10.435 2.290 12.235 2.460 ;
        RECT 10.435 2.050 10.685 2.290 ;
        RECT 10.855 1.950 11.895 2.120 ;
        RECT 10.855 1.880 11.025 1.950 ;
        RECT 9.030 1.540 9.350 1.800 ;
        RECT 9.735 1.710 11.025 1.880 ;
        RECT 11.195 1.540 11.395 1.780 ;
        RECT 9.030 1.470 10.395 1.540 ;
        RECT 9.180 1.370 10.395 1.470 ;
        RECT 7.145 1.130 9.010 1.300 ;
        RECT 10.065 1.225 10.395 1.370 ;
        RECT 10.995 1.210 11.395 1.540 ;
        RECT 6.665 0.765 6.930 1.095 ;
        RECT 9.495 0.960 9.825 1.200 ;
        RECT 11.565 1.040 11.895 1.950 ;
        RECT 7.100 0.790 9.825 0.960 ;
        RECT 9.995 0.870 11.895 1.040 ;
        RECT 7.100 0.545 7.270 0.790 ;
        RECT 9.995 0.620 10.165 0.870 ;
        RECT 12.065 0.700 12.235 2.290 ;
        RECT 1.165 0.255 3.390 0.425 ;
        RECT 3.575 0.085 4.065 0.360 ;
        RECT 4.805 0.085 5.165 0.360 ;
        RECT 6.325 0.255 7.270 0.545 ;
        RECT 7.890 0.085 8.220 0.620 ;
        RECT 9.190 0.290 10.165 0.620 ;
        RECT 10.730 0.085 11.200 0.680 ;
        RECT 11.690 0.450 12.235 0.700 ;
        RECT 12.440 1.685 12.795 2.980 ;
        RECT 12.975 1.820 13.305 3.245 ;
        RECT 12.440 1.355 12.810 1.685 ;
        RECT 12.440 0.350 12.795 1.355 ;
        RECT 12.975 0.085 13.305 1.130 ;
        RECT 0.000 -0.085 13.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 3.515 1.580 3.685 1.750 ;
        RECT 7.835 1.580 8.005 1.750 ;
        RECT 11.195 1.580 11.365 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
  END
END sky130_fd_sc_hs__sdfrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.260 4.640 1.590 ;
        RECT 3.965 1.180 4.195 1.260 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.810 2.100 1.265 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 3.935 2.105 4.225 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 10.655 2.105 10.945 2.150 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 3.935 1.920 4.225 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
        RECT 10.655 1.920 10.945 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.440 3.275 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.660 1.795 1.835 ;
        RECT 0.455 1.490 2.725 1.660 ;
        RECT 2.395 1.260 2.725 1.490 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.175 1.140 5.590 1.240 ;
        RECT 0.005 0.955 0.985 0.990 ;
        RECT 4.175 0.955 9.105 1.140 ;
        RECT 12.455 1.050 13.435 1.240 ;
        RECT 0.005 0.920 9.105 0.955 ;
        RECT 11.460 0.920 13.435 1.050 ;
        RECT 0.005 0.245 13.435 0.920 ;
        RECT 0.000 0.000 13.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.630 3.520 ;
        RECT 8.145 1.555 9.665 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.440 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 13.070 1.130 13.325 2.980 ;
        RECT 12.995 0.350 13.325 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.440 3.415 ;
        RECT 0.115 2.175 0.445 2.980 ;
        RECT 0.615 2.345 0.945 3.245 ;
        RECT 1.485 2.515 2.555 2.980 ;
        RECT 3.095 2.685 3.425 3.245 ;
        RECT 3.665 2.560 3.995 2.980 ;
        RECT 4.705 2.730 5.035 3.245 ;
        RECT 5.825 2.560 6.075 2.725 ;
        RECT 3.665 2.515 6.075 2.560 ;
        RECT 1.485 2.390 6.075 2.515 ;
        RECT 1.485 2.345 3.995 2.390 ;
        RECT 3.445 2.330 3.995 2.345 ;
        RECT 0.115 2.005 2.705 2.175 ;
        RECT 0.115 1.265 0.285 2.005 ;
        RECT 2.035 1.830 2.705 2.005 ;
        RECT 0.115 1.050 1.375 1.265 ;
        RECT 3.445 1.090 3.615 2.330 ;
        RECT 3.785 1.830 4.165 2.160 ;
        RECT 4.335 1.990 4.585 2.220 ;
        RECT 4.335 1.820 4.980 1.990 ;
        RECT 5.155 1.875 5.620 2.220 ;
        RECT 5.825 2.215 6.075 2.390 ;
        RECT 6.250 2.490 6.880 2.725 ;
        RECT 7.205 2.660 7.540 3.245 ;
        RECT 7.745 2.490 8.075 2.745 ;
        RECT 6.250 2.385 8.075 2.490 ;
        RECT 6.710 2.320 8.075 2.385 ;
        RECT 5.825 2.045 6.540 2.215 ;
        RECT 5.155 1.820 6.200 1.875 ;
        RECT 4.810 1.630 4.980 1.820 ;
        RECT 4.810 1.300 5.280 1.630 ;
        RECT 5.450 1.545 6.200 1.820 ;
        RECT 4.810 1.090 4.980 1.300 ;
        RECT 5.450 1.130 5.620 1.545 ;
        RECT 6.370 1.370 6.540 2.045 ;
        RECT 0.115 0.420 0.365 1.050 ;
        RECT 1.045 0.935 1.375 1.050 ;
        RECT 2.270 0.920 3.615 1.090 ;
        RECT 4.365 0.920 4.980 1.090 ;
        RECT 0.545 0.085 0.875 0.880 ;
        RECT 1.105 0.425 1.435 0.640 ;
        RECT 2.270 0.595 2.600 0.920 ;
        RECT 3.090 0.425 3.605 0.715 ;
        RECT 1.105 0.255 3.605 0.425 ;
        RECT 3.785 0.085 3.955 0.750 ;
        RECT 4.365 0.350 4.535 0.920 ;
        RECT 4.715 0.085 4.965 0.750 ;
        RECT 5.150 0.425 5.620 1.130 ;
        RECT 5.790 1.200 6.540 1.370 ;
        RECT 5.790 0.595 5.960 1.200 ;
        RECT 6.710 1.030 6.880 2.320 ;
        RECT 6.140 0.860 6.880 1.030 ;
        RECT 7.050 1.090 7.325 1.805 ;
        RECT 7.495 1.575 7.665 2.320 ;
        RECT 7.835 1.815 8.165 2.150 ;
        RECT 8.385 1.745 8.555 3.245 ;
        RECT 8.725 1.715 9.005 2.755 ;
        RECT 9.290 2.550 10.315 2.880 ;
        RECT 9.245 2.125 9.975 2.380 ;
        RECT 7.495 1.260 8.315 1.575 ;
        RECT 8.725 1.090 8.895 1.715 ;
        RECT 9.245 1.270 9.415 2.125 ;
        RECT 10.145 1.955 10.315 2.550 ;
        RECT 10.485 2.520 10.735 3.245 ;
        RECT 10.945 2.520 11.310 2.980 ;
        RECT 7.050 0.920 8.895 1.090 ;
        RECT 9.065 0.940 9.415 1.270 ;
        RECT 9.585 1.785 10.315 1.955 ;
        RECT 10.640 1.820 10.970 2.150 ;
        RECT 9.585 1.265 9.755 1.785 ;
        RECT 11.140 1.615 11.310 2.520 ;
        RECT 11.480 2.100 11.810 3.245 ;
        RECT 11.980 2.100 12.310 2.980 ;
        RECT 12.085 1.630 12.310 2.100 ;
        RECT 12.540 1.820 12.870 3.245 ;
        RECT 9.985 1.445 11.735 1.615 ;
        RECT 9.985 1.435 10.315 1.445 ;
        RECT 11.065 1.265 11.395 1.275 ;
        RECT 9.585 1.095 11.395 1.265 ;
        RECT 6.140 0.595 6.470 0.860 ;
        RECT 7.050 0.580 8.100 0.750 ;
        RECT 8.270 0.595 8.655 0.920 ;
        RECT 7.050 0.425 7.220 0.580 ;
        RECT 5.150 0.255 7.220 0.425 ;
        RECT 7.930 0.425 8.100 0.580 ;
        RECT 9.065 0.425 9.235 0.940 ;
        RECT 9.585 0.770 9.755 1.095 ;
        RECT 11.565 0.925 11.735 1.445 ;
        RECT 7.430 0.085 7.760 0.410 ;
        RECT 7.930 0.255 9.235 0.425 ;
        RECT 9.405 0.350 9.755 0.770 ;
        RECT 10.195 0.085 10.525 0.810 ;
        RECT 11.010 0.755 11.735 0.925 ;
        RECT 12.085 1.300 12.870 1.630 ;
        RECT 11.010 0.350 11.340 0.755 ;
        RECT 11.570 0.085 11.905 0.585 ;
        RECT 12.085 0.350 12.335 1.300 ;
        RECT 12.565 0.085 12.815 1.130 ;
        RECT 0.000 -0.085 13.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 10.715 1.950 10.885 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
  END
END sky130_fd_sc_hs__sdfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.400 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.260 4.645 1.590 ;
        RECT 3.965 1.180 4.195 1.260 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.810 2.100 1.265 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 3.935 2.105 4.225 2.150 ;
        RECT 8.255 2.105 8.545 2.150 ;
        RECT 11.135 2.105 11.425 2.150 ;
        RECT 3.935 1.965 11.425 2.105 ;
        RECT 3.935 1.920 4.225 1.965 ;
        RECT 8.255 1.920 8.545 1.965 ;
        RECT 11.135 1.920 11.425 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.480 3.275 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.660 1.795 1.835 ;
        RECT 0.605 1.490 2.705 1.660 ;
        RECT 2.375 1.260 2.705 1.490 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.200 0.955 9.500 1.240 ;
        RECT 12.985 1.140 14.395 1.240 ;
        RECT 0.995 0.920 9.500 0.955 ;
        RECT 11.995 0.920 14.395 1.140 ;
        RECT 0.005 0.245 14.395 0.920 ;
        RECT 0.000 0.000 14.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.590 3.520 ;
        RECT 8.120 1.555 9.780 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.400 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 13.525 1.410 13.785 2.980 ;
        RECT 13.525 0.350 13.855 1.410 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.400 3.415 ;
        RECT 0.115 2.175 0.445 2.980 ;
        RECT 0.615 2.345 1.565 3.245 ;
        RECT 2.105 2.515 2.435 2.980 ;
        RECT 3.095 2.685 3.425 3.245 ;
        RECT 3.615 2.560 3.995 2.980 ;
        RECT 4.705 2.730 5.035 3.245 ;
        RECT 5.745 2.560 5.995 2.725 ;
        RECT 3.615 2.515 5.995 2.560 ;
        RECT 2.105 2.390 5.995 2.515 ;
        RECT 6.195 2.490 6.870 2.725 ;
        RECT 7.150 2.660 7.485 3.245 ;
        RECT 7.690 2.490 8.020 2.725 ;
        RECT 6.195 2.475 8.020 2.490 ;
        RECT 2.105 2.345 3.995 2.390 ;
        RECT 3.445 2.330 3.995 2.345 ;
        RECT 0.115 2.005 2.705 2.175 ;
        RECT 0.115 1.265 0.285 2.005 ;
        RECT 2.375 1.830 2.705 2.005 ;
        RECT 3.445 1.310 3.615 2.330 ;
        RECT 5.745 2.305 5.995 2.390 ;
        RECT 6.700 2.320 8.020 2.475 ;
        RECT 8.250 2.320 8.580 3.245 ;
        RECT 3.785 1.830 4.165 2.160 ;
        RECT 4.335 1.990 4.585 2.220 ;
        RECT 4.335 1.820 4.985 1.990 ;
        RECT 0.115 0.935 1.140 1.265 ;
        RECT 2.875 1.140 3.615 1.310 ;
        RECT 4.815 1.625 4.985 1.820 ;
        RECT 5.155 1.965 5.485 2.220 ;
        RECT 5.745 2.135 6.530 2.305 ;
        RECT 5.155 1.795 6.190 1.965 ;
        RECT 5.475 1.635 6.190 1.795 ;
        RECT 4.815 1.295 5.305 1.625 ;
        RECT 0.115 0.350 0.365 0.935 ;
        RECT 2.875 0.845 3.045 1.140 ;
        RECT 4.815 1.090 4.985 1.295 ;
        RECT 5.475 1.125 5.645 1.635 ;
        RECT 6.360 1.465 6.530 2.135 ;
        RECT 4.390 0.920 4.985 1.090 ;
        RECT 0.545 0.085 0.875 0.765 ;
        RECT 1.105 0.425 1.435 0.640 ;
        RECT 2.270 0.595 3.045 0.845 ;
        RECT 3.215 0.425 3.545 0.845 ;
        RECT 1.105 0.255 3.545 0.425 ;
        RECT 3.715 0.085 4.045 0.845 ;
        RECT 4.390 0.350 4.560 0.920 ;
        RECT 4.740 0.085 5.070 0.750 ;
        RECT 5.240 0.500 5.645 1.125 ;
        RECT 5.815 1.295 6.530 1.465 ;
        RECT 5.815 0.670 6.145 1.295 ;
        RECT 6.700 1.125 6.870 2.320 ;
        RECT 6.315 0.955 6.870 1.125 ;
        RECT 7.040 1.090 7.315 2.075 ;
        RECT 7.485 1.575 7.655 2.320 ;
        RECT 7.825 1.795 8.515 2.150 ;
        RECT 8.750 1.715 9.115 2.755 ;
        RECT 9.320 2.520 10.390 2.850 ;
        RECT 10.560 2.730 11.240 3.245 ;
        RECT 11.410 2.560 11.740 2.980 ;
        RECT 9.320 1.840 9.600 2.520 ;
        RECT 7.485 1.260 8.420 1.575 ;
        RECT 8.750 1.130 8.920 1.715 ;
        RECT 9.785 1.335 10.050 2.330 ;
        RECT 8.590 1.090 8.920 1.130 ;
        RECT 6.315 0.670 6.645 0.955 ;
        RECT 7.040 0.920 8.920 1.090 ;
        RECT 7.040 0.580 8.420 0.750 ;
        RECT 8.590 0.595 8.920 0.920 ;
        RECT 9.090 1.005 10.050 1.335 ;
        RECT 10.220 1.200 10.390 2.520 ;
        RECT 10.560 2.390 11.740 2.560 ;
        RECT 10.560 1.750 10.850 2.390 ;
        RECT 11.110 1.920 11.440 2.220 ;
        RECT 11.945 1.940 12.275 3.245 ;
        RECT 12.445 1.940 12.775 2.980 ;
        RECT 10.560 1.580 12.230 1.750 ;
        RECT 10.560 1.370 10.850 1.580 ;
        RECT 11.020 1.200 11.890 1.410 ;
        RECT 10.220 1.110 11.890 1.200 ;
        RECT 10.220 1.030 11.190 1.110 ;
        RECT 7.040 0.500 7.210 0.580 ;
        RECT 5.240 0.330 7.210 0.500 ;
        RECT 8.250 0.425 8.420 0.580 ;
        RECT 9.090 0.425 9.260 1.005 ;
        RECT 10.220 0.810 10.390 1.030 ;
        RECT 12.060 0.940 12.230 1.580 ;
        RECT 9.430 0.480 10.390 0.810 ;
        RECT 7.605 0.085 8.080 0.410 ;
        RECT 8.250 0.255 9.260 0.425 ;
        RECT 10.755 0.085 11.085 0.810 ;
        RECT 11.545 0.770 12.230 0.940 ;
        RECT 12.605 1.630 12.775 1.940 ;
        RECT 13.005 1.820 13.335 3.245 ;
        RECT 13.955 1.820 14.285 3.245 ;
        RECT 12.605 1.300 13.355 1.630 ;
        RECT 11.545 0.350 11.875 0.770 ;
        RECT 12.105 0.085 12.435 0.600 ;
        RECT 12.605 0.350 12.865 1.300 ;
        RECT 13.095 0.085 13.345 1.130 ;
        RECT 14.035 0.085 14.285 1.130 ;
        RECT 0.000 -0.085 14.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 8.315 1.950 8.485 2.120 ;
        RECT 11.195 1.950 11.365 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
  END
END sky130_fd_sc_hs__sdfrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.880 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.260 4.635 1.590 ;
        RECT 3.965 1.180 4.195 1.260 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.810 2.100 1.265 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.411000 ;
    PORT
      LAYER met1 ;
        RECT 3.935 2.105 4.225 2.150 ;
        RECT 7.775 2.105 8.065 2.150 ;
        RECT 10.655 2.105 10.945 2.150 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 3.935 1.920 4.225 1.965 ;
        RECT 7.775 1.920 8.065 1.965 ;
        RECT 10.655 1.920 10.945 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.440 3.275 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.660 1.795 1.835 ;
        RECT 0.605 1.490 2.735 1.660 ;
        RECT 2.405 1.260 2.735 1.490 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.175 1.140 8.630 1.240 ;
        RECT 4.175 0.955 9.105 1.140 ;
        RECT 0.995 0.920 9.105 0.955 ;
        RECT 11.565 0.920 14.875 1.240 ;
        RECT 0.005 0.245 14.875 0.920 ;
        RECT 0.000 0.000 14.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 15.070 3.520 ;
        RECT 8.125 1.555 9.645 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.880 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 13.085 1.940 13.415 2.980 ;
        RECT 14.065 1.940 14.280 2.980 ;
        RECT 13.085 1.770 14.755 1.940 ;
        RECT 14.085 1.300 14.755 1.770 ;
        RECT 14.085 1.100 14.255 1.300 ;
        RECT 12.535 0.930 14.255 1.100 ;
        RECT 12.535 0.350 12.865 0.930 ;
        RECT 14.085 0.350 14.255 0.930 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.880 3.415 ;
        RECT 0.115 2.175 0.445 2.980 ;
        RECT 0.615 2.345 1.565 3.245 ;
        RECT 2.105 2.515 2.435 2.980 ;
        RECT 3.095 2.685 3.425 3.245 ;
        RECT 3.615 2.560 3.995 2.980 ;
        RECT 4.705 2.730 5.035 3.245 ;
        RECT 5.745 2.560 6.075 2.755 ;
        RECT 3.615 2.515 6.075 2.560 ;
        RECT 2.105 2.390 6.075 2.515 ;
        RECT 6.245 2.490 6.885 2.755 ;
        RECT 7.170 2.660 7.520 3.245 ;
        RECT 7.725 2.490 8.055 2.755 ;
        RECT 6.245 2.425 8.055 2.490 ;
        RECT 2.105 2.345 3.995 2.390 ;
        RECT 3.445 2.330 3.995 2.345 ;
        RECT 0.115 2.005 2.705 2.175 ;
        RECT 0.115 1.265 0.285 2.005 ;
        RECT 2.375 1.830 2.705 2.005 ;
        RECT 0.115 0.935 1.140 1.265 ;
        RECT 3.445 1.090 3.615 2.330 ;
        RECT 5.745 2.255 6.075 2.390 ;
        RECT 6.715 2.320 8.055 2.425 ;
        RECT 3.785 1.830 4.165 2.160 ;
        RECT 4.335 1.990 4.585 2.220 ;
        RECT 4.335 1.820 4.975 1.990 ;
        RECT 4.805 1.575 4.975 1.820 ;
        RECT 5.155 1.915 5.485 2.220 ;
        RECT 5.745 2.085 6.545 2.255 ;
        RECT 5.155 1.745 6.205 1.915 ;
        RECT 5.450 1.585 6.205 1.745 ;
        RECT 4.805 1.245 5.280 1.575 ;
        RECT 4.805 1.090 4.975 1.245 ;
        RECT 0.115 0.350 0.365 0.935 ;
        RECT 2.565 0.920 3.615 1.090 ;
        RECT 4.365 0.920 4.975 1.090 ;
        RECT 5.450 1.075 5.620 1.585 ;
        RECT 6.375 1.415 6.545 2.085 ;
        RECT 2.565 0.845 2.735 0.920 ;
        RECT 0.545 0.085 0.875 0.765 ;
        RECT 1.105 0.425 1.435 0.640 ;
        RECT 2.270 0.595 2.735 0.845 ;
        RECT 3.225 0.425 3.555 0.750 ;
        RECT 1.105 0.255 3.555 0.425 ;
        RECT 3.725 0.085 4.055 0.750 ;
        RECT 4.365 0.350 4.535 0.920 ;
        RECT 4.715 0.085 4.965 0.750 ;
        RECT 5.145 0.500 5.620 1.075 ;
        RECT 5.790 1.245 6.545 1.415 ;
        RECT 5.790 0.670 5.960 1.245 ;
        RECT 6.715 1.075 6.885 2.320 ;
        RECT 6.140 0.905 6.885 1.075 ;
        RECT 7.055 1.090 7.325 1.945 ;
        RECT 7.495 1.575 7.665 2.320 ;
        RECT 7.835 1.820 8.145 2.150 ;
        RECT 8.365 1.745 8.535 3.245 ;
        RECT 8.735 1.575 9.065 2.755 ;
        RECT 9.270 2.550 10.295 2.880 ;
        RECT 7.495 1.260 8.315 1.575 ;
        RECT 8.485 1.405 9.065 1.575 ;
        RECT 9.245 2.065 9.955 2.380 ;
        RECT 8.485 1.090 8.655 1.405 ;
        RECT 9.245 1.235 9.415 2.065 ;
        RECT 10.125 1.895 10.295 2.550 ;
        RECT 10.465 2.520 10.795 3.245 ;
        RECT 11.000 2.520 11.330 2.980 ;
        RECT 7.055 0.920 8.655 1.090 ;
        RECT 6.140 0.670 6.470 0.905 ;
        RECT 7.055 0.580 8.100 0.750 ;
        RECT 8.270 0.595 8.655 0.920 ;
        RECT 8.825 0.905 9.415 1.235 ;
        RECT 9.585 1.725 10.295 1.895 ;
        RECT 10.585 1.820 10.915 2.150 ;
        RECT 9.585 1.055 9.755 1.725 ;
        RECT 11.160 1.555 11.330 2.520 ;
        RECT 11.650 1.820 11.900 3.245 ;
        RECT 12.100 1.600 12.430 2.700 ;
        RECT 12.635 1.820 12.885 3.245 ;
        RECT 13.615 2.110 13.865 3.245 ;
        RECT 14.470 2.110 14.765 3.245 ;
        RECT 10.015 1.385 11.585 1.555 ;
        RECT 10.015 1.225 10.345 1.385 ;
        RECT 10.915 1.055 11.245 1.215 ;
        RECT 7.055 0.500 7.225 0.580 ;
        RECT 5.145 0.330 7.225 0.500 ;
        RECT 7.930 0.425 8.100 0.580 ;
        RECT 8.825 0.425 8.995 0.905 ;
        RECT 9.585 0.885 11.245 1.055 ;
        RECT 9.585 0.735 9.755 0.885 ;
        RECT 7.430 0.085 7.760 0.410 ;
        RECT 7.930 0.255 8.995 0.425 ;
        RECT 9.165 0.405 9.755 0.735 ;
        RECT 11.415 0.715 11.585 1.385 ;
        RECT 10.140 0.085 10.580 0.680 ;
        RECT 11.040 0.385 11.585 0.715 ;
        RECT 11.755 1.270 13.850 1.600 ;
        RECT 11.755 0.350 11.925 1.270 ;
        RECT 12.105 0.085 12.365 1.100 ;
        RECT 13.035 0.085 13.905 0.760 ;
        RECT 14.435 0.085 14.765 1.130 ;
        RECT 0.000 -0.085 14.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 3.995 1.950 4.165 2.120 ;
        RECT 7.835 1.950 8.005 2.120 ;
        RECT 10.715 1.950 10.885 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
  END
END sky130_fd_sc_hs__sdfrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.400 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.275 1.180 3.715 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.790 1.585 2.120 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.140 2.765 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.620 0.835 1.850 ;
        RECT 0.505 1.450 2.045 1.620 ;
        RECT 1.795 1.260 2.045 1.450 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.735 7.585 1.780 ;
        RECT 9.695 1.735 9.985 1.780 ;
        RECT 7.295 1.595 9.985 1.735 ;
        RECT 7.295 1.550 7.585 1.595 ;
        RECT 9.695 1.550 9.985 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.400 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.840 1.035 4.320 1.240 ;
        RECT 2.840 0.920 4.880 1.035 ;
        RECT 7.390 0.920 9.225 1.140 ;
        RECT 11.515 0.920 14.395 1.240 ;
        RECT 0.005 0.245 14.395 0.920 ;
        RECT 0.000 0.000 14.400 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.590 3.520 ;
        RECT 7.405 1.555 8.470 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.400 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.535700 ;
    PORT
      LAYER li1 ;
        RECT 13.955 0.350 14.290 2.980 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.535700 ;
    PORT
      LAYER li1 ;
        RECT 12.450 1.820 12.705 2.980 ;
        RECT 12.450 1.130 12.620 1.820 ;
        RECT 12.125 0.350 12.620 1.130 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.400 3.415 ;
        RECT 0.115 2.460 0.365 2.980 ;
        RECT 0.565 2.630 0.895 3.245 ;
        RECT 1.435 2.800 1.945 2.960 ;
        RECT 1.435 2.630 2.385 2.800 ;
        RECT 2.555 2.660 2.820 3.245 ;
        RECT 3.575 2.660 3.905 3.245 ;
        RECT 4.105 2.905 5.810 3.075 ;
        RECT 2.215 2.490 2.385 2.630 ;
        RECT 4.105 2.550 4.355 2.905 ;
        RECT 0.115 2.290 2.045 2.460 ;
        RECT 0.115 1.280 0.335 2.290 ;
        RECT 1.795 1.830 2.045 2.290 ;
        RECT 2.215 2.380 3.795 2.490 ;
        RECT 4.590 2.380 4.925 2.735 ;
        RECT 2.215 2.320 4.925 2.380 ;
        RECT 5.120 2.370 5.450 2.735 ;
        RECT 0.115 0.950 1.140 1.280 ;
        RECT 2.215 1.090 2.385 2.320 ;
        RECT 3.625 2.210 4.925 2.320 ;
        RECT 0.115 0.350 0.445 0.950 ;
        RECT 1.505 0.920 2.385 1.090 ;
        RECT 2.935 1.990 3.455 2.150 ;
        RECT 2.935 1.820 4.215 1.990 ;
        RECT 2.935 1.010 3.105 1.820 ;
        RECT 3.885 1.220 4.215 1.820 ;
        RECT 0.615 0.085 0.945 0.780 ;
        RECT 1.505 0.350 1.835 0.920 ;
        RECT 2.325 0.085 2.655 0.750 ;
        RECT 2.935 0.340 3.200 1.010 ;
        RECT 3.380 0.085 3.710 1.010 ;
        RECT 3.880 0.425 4.210 1.010 ;
        RECT 4.420 0.925 4.590 2.210 ;
        RECT 4.760 1.370 5.030 2.040 ;
        RECT 4.420 0.595 4.690 0.925 ;
        RECT 4.860 0.425 5.030 1.370 ;
        RECT 3.880 0.255 5.030 0.425 ;
        RECT 5.200 1.520 5.370 2.370 ;
        RECT 5.640 2.255 5.810 2.905 ;
        RECT 6.175 2.425 6.425 3.245 ;
        RECT 6.595 2.905 7.445 3.075 ;
        RECT 6.595 2.255 6.765 2.905 ;
        RECT 5.640 2.085 6.765 2.255 ;
        RECT 5.640 2.020 5.810 2.085 ;
        RECT 5.540 1.690 5.810 2.020 ;
        RECT 6.935 1.915 7.105 2.735 ;
        RECT 7.275 2.120 7.445 2.905 ;
        RECT 7.615 2.295 7.785 3.245 ;
        RECT 8.530 2.905 10.380 3.075 ;
        RECT 7.985 2.520 8.315 2.755 ;
        RECT 8.530 2.690 8.860 2.905 ;
        RECT 9.580 2.520 9.830 2.735 ;
        RECT 10.050 2.520 10.380 2.905 ;
        RECT 10.580 2.520 10.750 3.245 ;
        RECT 10.950 2.520 11.280 2.980 ;
        RECT 7.985 2.350 9.830 2.520 ;
        RECT 7.985 2.290 8.315 2.350 ;
        RECT 9.580 2.290 9.830 2.350 ;
        RECT 11.110 2.265 11.280 2.520 ;
        RECT 9.045 2.120 9.380 2.180 ;
        RECT 10.000 2.120 11.280 2.265 ;
        RECT 11.500 2.350 11.750 2.980 ;
        RECT 11.950 2.520 12.280 3.245 ;
        RECT 11.500 2.180 12.235 2.350 ;
        RECT 7.275 1.950 8.830 2.120 ;
        RECT 6.050 1.690 7.105 1.915 ;
        RECT 5.200 1.350 7.110 1.520 ;
        RECT 5.200 0.350 5.450 1.350 ;
        RECT 6.725 1.190 7.110 1.350 ;
        RECT 7.295 1.245 7.625 1.780 ;
        RECT 8.660 1.680 8.830 1.950 ;
        RECT 9.045 2.095 11.280 2.120 ;
        RECT 9.045 1.950 10.170 2.095 ;
        RECT 11.110 1.970 11.280 2.095 ;
        RECT 9.045 1.850 9.380 1.950 ;
        RECT 5.815 0.905 6.485 1.180 ;
        RECT 6.940 1.075 7.110 1.190 ;
        RECT 7.835 1.075 8.165 1.450 ;
        RECT 8.660 1.350 8.990 1.680 ;
        RECT 6.940 0.905 8.165 1.075 ;
        RECT 9.210 1.050 9.380 1.850 ;
        RECT 10.585 1.780 10.915 1.925 ;
        RECT 9.725 1.550 10.915 1.780 ;
        RECT 11.110 1.640 11.895 1.970 ;
        RECT 10.585 1.255 10.915 1.550 ;
        RECT 12.065 1.470 12.235 2.180 ;
        RECT 11.225 1.300 12.235 1.470 ;
        RECT 13.005 1.550 13.255 2.875 ;
        RECT 13.455 1.995 13.785 3.245 ;
        RECT 5.815 0.735 6.770 0.905 ;
        RECT 6.020 0.085 6.370 0.565 ;
        RECT 6.600 0.350 6.930 0.735 ;
        RECT 7.500 0.085 8.295 0.735 ;
        RECT 8.785 0.350 9.380 1.050 ;
        RECT 9.620 1.070 9.950 1.230 ;
        RECT 11.225 1.070 11.395 1.300 ;
        RECT 13.005 1.220 13.785 1.550 ;
        RECT 13.005 1.130 13.255 1.220 ;
        RECT 9.620 0.900 11.395 1.070 ;
        RECT 10.285 0.085 10.895 0.680 ;
        RECT 11.065 0.350 11.395 0.900 ;
        RECT 11.625 0.085 11.955 1.130 ;
        RECT 12.840 0.540 13.255 1.130 ;
        RECT 13.455 0.085 13.785 1.050 ;
        RECT 0.000 -0.085 14.400 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 7.355 1.580 7.525 1.750 ;
        RECT 9.755 1.580 9.925 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
  END
END sky130_fd_sc_hs__sdfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfsbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.760 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.715 1.180 4.195 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.385 0.440 1.795 1.230 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.805 0.950 3.205 1.620 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.570 1.085 1.800 ;
        RECT 0.425 1.400 2.295 1.570 ;
        RECT 1.965 0.900 2.295 1.400 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.735 8.065 1.780 ;
        RECT 13.055 1.735 13.345 1.780 ;
        RECT 7.775 1.595 13.345 1.735 ;
        RECT 7.775 1.550 8.065 1.595 ;
        RECT 13.055 1.550 13.345 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 17.760 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.290 0.955 4.770 1.240 ;
        RECT 3.290 0.920 7.260 0.955 ;
        RECT 8.840 0.920 11.320 1.140 ;
        RECT 14.240 0.920 17.755 1.240 ;
        RECT 0.005 0.245 17.755 0.920 ;
        RECT 0.000 0.000 17.760 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 17.950 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 17.760 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 16.865 1.820 17.225 2.980 ;
        RECT 17.055 1.130 17.225 1.820 ;
        RECT 16.885 0.350 17.225 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 14.850 1.410 15.105 2.980 ;
        RECT 14.850 0.350 15.235 1.410 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 17.760 3.415 ;
        RECT 0.085 2.140 0.465 2.980 ;
        RECT 0.635 2.310 0.965 3.245 ;
        RECT 1.505 2.480 1.955 2.980 ;
        RECT 2.495 2.650 2.845 3.245 ;
        RECT 3.525 2.650 4.220 3.245 ;
        RECT 4.390 2.905 6.240 3.075 ;
        RECT 1.505 2.310 3.885 2.480 ;
        RECT 4.390 2.470 4.720 2.905 ;
        RECT 0.085 1.970 2.105 2.140 ;
        RECT 0.085 1.230 0.255 1.970 ;
        RECT 1.775 1.810 2.105 1.970 ;
        RECT 0.085 0.900 1.145 1.230 ;
        RECT 0.085 0.350 0.445 0.900 ;
        RECT 2.465 0.730 2.635 2.310 ;
        RECT 3.715 2.300 3.885 2.310 ;
        RECT 4.890 2.300 5.370 2.735 ;
        RECT 3.075 1.960 3.545 2.140 ;
        RECT 3.715 2.130 5.370 2.300 ;
        RECT 5.540 2.295 5.900 2.735 ;
        RECT 3.075 1.790 4.720 1.960 ;
        RECT 3.375 1.010 3.545 1.790 ;
        RECT 4.390 1.350 4.720 1.790 ;
        RECT 0.615 0.085 1.020 0.680 ;
        RECT 1.965 0.560 2.635 0.730 ;
        RECT 1.965 0.400 2.350 0.560 ;
        RECT 2.840 0.085 3.170 0.780 ;
        RECT 3.375 0.340 3.650 1.010 ;
        RECT 3.830 0.085 4.160 1.010 ;
        RECT 4.330 0.425 4.660 1.010 ;
        RECT 4.890 0.845 5.060 2.130 ;
        RECT 5.230 1.290 5.560 1.960 ;
        RECT 4.890 0.595 5.220 0.845 ;
        RECT 5.390 0.425 5.560 1.290 ;
        RECT 5.730 0.800 5.900 2.295 ;
        RECT 6.070 2.335 6.240 2.905 ;
        RECT 6.410 2.505 6.985 3.245 ;
        RECT 7.155 2.905 8.165 3.075 ;
        RECT 7.155 2.335 7.325 2.905 ;
        RECT 6.070 2.165 7.325 2.335 ;
        RECT 7.495 2.295 7.825 2.735 ;
        RECT 6.070 0.970 6.305 2.165 ;
        RECT 7.495 1.995 7.665 2.295 ;
        RECT 7.995 2.220 8.165 2.905 ;
        RECT 8.335 2.390 8.665 3.245 ;
        RECT 8.925 2.300 9.255 2.980 ;
        RECT 9.425 2.470 9.675 3.245 ;
        RECT 9.875 2.905 11.105 3.075 ;
        RECT 9.875 2.300 10.125 2.905 ;
        RECT 7.995 2.050 8.565 2.220 ;
        RECT 8.925 2.130 10.125 2.300 ;
        RECT 9.875 2.100 10.125 2.130 ;
        RECT 10.325 2.210 10.575 2.700 ;
        RECT 10.775 2.380 11.105 2.905 ;
        RECT 11.365 2.885 12.740 3.055 ;
        RECT 11.365 2.385 11.620 2.885 ;
        RECT 11.820 2.310 12.220 2.715 ;
        RECT 12.410 2.520 12.740 2.885 ;
        RECT 12.940 2.520 13.110 3.245 ;
        RECT 13.310 2.310 13.640 2.980 ;
        RECT 13.870 2.480 14.315 2.910 ;
        RECT 11.820 2.210 13.975 2.310 ;
        RECT 10.325 2.140 13.975 2.210 ;
        RECT 6.635 1.735 7.665 1.995 ;
        RECT 6.475 1.395 7.665 1.565 ;
        RECT 7.835 1.550 8.225 1.880 ;
        RECT 6.475 0.800 6.645 1.395 ;
        RECT 7.355 1.380 7.665 1.395 ;
        RECT 8.395 1.515 8.565 2.050 ;
        RECT 10.325 2.040 12.390 2.140 ;
        RECT 8.735 1.870 9.065 1.960 ;
        RECT 8.735 1.700 12.050 1.870 ;
        RECT 8.735 1.685 9.065 1.700 ;
        RECT 10.380 1.515 11.390 1.530 ;
        RECT 6.815 1.040 7.145 1.225 ;
        RECT 7.355 1.210 8.050 1.380 ;
        RECT 8.395 1.345 11.390 1.515 ;
        RECT 7.880 1.175 8.050 1.210 ;
        RECT 10.380 1.200 11.390 1.345 ;
        RECT 6.815 0.870 7.710 1.040 ;
        RECT 7.880 0.900 8.860 1.175 ;
        RECT 9.030 1.005 10.210 1.175 ;
        RECT 5.730 0.470 6.645 0.800 ;
        RECT 4.330 0.255 5.560 0.425 ;
        RECT 6.815 0.085 7.150 0.700 ;
        RECT 7.380 0.350 7.710 0.870 ;
        RECT 8.200 0.085 8.530 0.680 ;
        RECT 9.030 0.350 9.280 1.005 ;
        RECT 9.450 0.085 9.780 0.835 ;
        RECT 9.960 0.425 10.210 1.005 ;
        RECT 10.380 0.860 11.550 1.030 ;
        RECT 11.720 0.900 12.050 1.700 ;
        RECT 10.380 0.595 10.710 0.860 ;
        RECT 11.380 0.730 11.550 0.860 ;
        RECT 12.220 0.730 12.390 2.040 ;
        RECT 12.565 1.130 12.895 1.960 ;
        RECT 13.085 1.300 13.435 1.970 ;
        RECT 13.645 1.300 13.975 2.140 ;
        RECT 14.145 1.130 14.315 2.480 ;
        RECT 14.485 1.820 14.655 3.245 ;
        RECT 15.305 1.820 15.635 3.245 ;
        RECT 15.865 1.630 16.195 2.860 ;
        RECT 16.415 1.820 16.665 3.245 ;
        RECT 17.395 1.820 17.645 3.245 ;
        RECT 15.865 1.300 16.885 1.630 ;
        RECT 12.565 0.960 14.315 1.130 ;
        RECT 10.880 0.425 11.210 0.690 ;
        RECT 9.960 0.255 11.210 0.425 ;
        RECT 11.380 0.400 12.390 0.730 ;
        RECT 13.260 0.085 13.590 0.790 ;
        RECT 13.770 0.350 14.100 0.960 ;
        RECT 14.350 0.085 14.680 0.790 ;
        RECT 15.405 0.085 15.655 1.130 ;
        RECT 15.865 0.450 16.220 1.300 ;
        RECT 16.455 0.085 16.705 1.130 ;
        RECT 17.395 0.085 17.645 1.130 ;
        RECT 0.000 -0.085 17.760 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 16.955 3.245 17.125 3.415 ;
        RECT 17.435 3.245 17.605 3.415 ;
        RECT 7.835 1.580 8.005 1.750 ;
        RECT 13.115 1.580 13.285 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
        RECT 17.435 -0.085 17.605 0.085 ;
  END
END sky130_fd_sc_hs__sdfsbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.180 3.715 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.820 1.580 2.150 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.140 2.805 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.610 0.835 1.950 ;
        RECT 0.425 1.440 2.045 1.610 ;
        RECT 0.425 1.280 0.680 1.440 ;
        RECT 1.790 1.260 2.045 1.440 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.735 7.585 1.780 ;
        RECT 10.655 1.735 10.945 1.780 ;
        RECT 7.295 1.595 10.945 1.735 ;
        RECT 7.295 1.550 7.585 1.595 ;
        RECT 10.655 1.550 10.945 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.920 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.865 0.955 4.415 1.240 ;
        RECT 6.565 0.955 9.455 1.140 ;
        RECT 2.865 0.920 9.455 0.955 ;
        RECT 11.845 0.920 13.820 1.240 ;
        RECT 0.085 0.245 13.820 0.920 ;
        RECT 0.000 0.000 13.920 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 14.110 3.520 ;
        RECT 7.455 1.525 8.515 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.920 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 13.565 1.050 13.815 2.980 ;
        RECT 13.380 0.350 13.815 1.050 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.920 3.415 ;
        RECT 0.085 2.490 0.360 2.980 ;
        RECT 0.560 2.660 0.890 3.245 ;
        RECT 1.430 2.660 2.385 2.910 ;
        RECT 2.565 2.830 2.895 3.245 ;
        RECT 2.215 2.490 3.405 2.660 ;
        RECT 3.575 2.580 3.905 3.245 ;
        RECT 4.105 2.895 5.845 3.065 ;
        RECT 4.105 2.580 4.275 2.895 ;
        RECT 0.085 2.320 2.045 2.490 ;
        RECT 0.085 2.300 0.360 2.320 ;
        RECT 0.085 1.110 0.255 2.300 ;
        RECT 1.790 1.830 2.045 2.320 ;
        RECT 0.890 1.110 1.220 1.270 ;
        RECT 0.085 0.940 1.220 1.110 ;
        RECT 2.215 1.090 2.385 2.490 ;
        RECT 3.235 2.410 3.405 2.490 ;
        RECT 4.445 2.410 5.005 2.725 ;
        RECT 3.235 2.240 5.005 2.410 ;
        RECT 5.175 2.265 5.505 2.725 ;
        RECT 5.675 2.515 5.845 2.895 ;
        RECT 6.225 2.685 6.475 3.245 ;
        RECT 6.645 2.895 7.495 3.065 ;
        RECT 6.645 2.515 6.815 2.895 ;
        RECT 5.675 2.345 6.815 2.515 ;
        RECT 0.085 0.350 0.525 0.940 ;
        RECT 1.555 0.920 2.385 1.090 ;
        RECT 2.975 1.820 4.215 2.070 ;
        RECT 2.975 1.010 3.145 1.820 ;
        RECT 3.885 1.350 4.215 1.820 ;
        RECT 0.695 0.085 1.025 0.770 ;
        RECT 1.555 0.350 1.885 0.920 ;
        RECT 2.375 0.085 2.705 0.750 ;
        RECT 2.975 0.350 3.305 1.010 ;
        RECT 3.475 0.085 3.805 1.010 ;
        RECT 3.975 0.425 4.225 1.130 ;
        RECT 4.445 0.765 4.615 2.240 ;
        RECT 4.785 1.105 5.005 2.070 ;
        RECT 5.175 1.445 5.345 2.265 ;
        RECT 5.675 1.945 5.845 2.345 ;
        RECT 6.985 2.175 7.155 2.725 ;
        RECT 5.515 1.775 5.845 1.945 ;
        RECT 6.015 2.005 7.155 2.175 ;
        RECT 7.325 2.140 7.495 2.895 ;
        RECT 7.665 2.310 7.915 3.245 ;
        RECT 8.585 2.905 10.430 3.075 ;
        RECT 8.115 2.520 8.365 2.725 ;
        RECT 8.585 2.690 8.915 2.905 ;
        RECT 9.565 2.520 9.895 2.735 ;
        RECT 10.100 2.560 10.430 2.905 ;
        RECT 10.630 2.560 10.800 3.245 ;
        RECT 8.115 2.350 9.895 2.520 ;
        RECT 11.000 2.390 11.370 2.980 ;
        RECT 6.015 1.795 6.345 2.005 ;
        RECT 7.325 1.970 7.945 2.140 ;
        RECT 5.515 1.615 5.730 1.775 ;
        RECT 6.650 1.605 6.935 1.835 ;
        RECT 5.900 1.445 6.935 1.605 ;
        RECT 7.145 1.540 7.555 1.800 ;
        RECT 7.775 1.750 7.945 1.970 ;
        RECT 8.115 1.920 8.365 2.350 ;
        RECT 9.090 1.790 9.365 2.180 ;
        RECT 9.565 1.960 9.895 2.350 ;
        RECT 10.065 2.220 11.370 2.390 ;
        RECT 11.540 2.390 11.870 2.980 ;
        RECT 12.070 2.560 12.320 3.245 ;
        RECT 11.540 2.220 11.940 2.390 ;
        RECT 10.065 1.790 10.235 2.220 ;
        RECT 11.200 2.050 11.370 2.220 ;
        RECT 7.775 1.580 8.840 1.750 ;
        RECT 9.090 1.620 10.235 1.790 ;
        RECT 5.175 1.435 6.935 1.445 ;
        RECT 5.175 1.275 6.070 1.435 ;
        RECT 6.650 1.370 6.935 1.435 ;
        RECT 8.670 1.450 8.840 1.580 ;
        RECT 7.760 1.370 8.430 1.410 ;
        RECT 4.785 0.935 5.205 1.105 ;
        RECT 4.445 0.595 4.865 0.765 ;
        RECT 5.035 0.425 5.205 0.935 ;
        RECT 3.975 0.255 5.205 0.425 ;
        RECT 5.375 0.385 5.625 1.275 ;
        RECT 6.240 1.030 6.480 1.265 ;
        RECT 6.650 1.200 8.430 1.370 ;
        RECT 7.760 1.120 8.430 1.200 ;
        RECT 8.670 1.120 9.000 1.450 ;
        RECT 6.240 0.860 7.005 1.030 ;
        RECT 9.195 0.940 9.365 1.620 ;
        RECT 10.685 1.380 11.030 2.050 ;
        RECT 11.200 1.380 11.600 2.050 ;
        RECT 9.790 1.210 10.460 1.310 ;
        RECT 11.770 1.210 11.940 2.220 ;
        RECT 9.790 1.040 11.940 1.210 ;
        RECT 12.530 1.995 12.860 2.875 ;
        RECT 13.030 1.995 13.360 3.245 ;
        RECT 12.530 1.550 12.700 1.995 ;
        RECT 12.530 1.220 13.395 1.550 ;
        RECT 9.790 0.980 11.770 1.040 ;
        RECT 12.530 1.005 12.700 1.220 ;
        RECT 6.115 0.085 6.445 0.690 ;
        RECT 6.675 0.570 7.005 0.860 ;
        RECT 7.455 0.085 8.305 0.940 ;
        RECT 8.795 0.350 9.365 0.940 ;
        RECT 10.825 0.085 11.155 0.810 ;
        RECT 11.395 0.350 11.770 0.980 ;
        RECT 12.370 0.870 12.700 1.005 ;
        RECT 11.955 0.540 12.700 0.870 ;
        RECT 12.880 0.085 13.210 1.050 ;
        RECT 0.000 -0.085 13.920 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 7.355 1.580 7.525 1.750 ;
        RECT 10.715 1.580 10.885 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
  END
END sky130_fd_sc_hs__sdfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfstp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.300 1.180 3.715 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.820 1.585 2.150 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.140 2.780 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.475 1.580 0.805 2.140 ;
        RECT 0.475 1.410 2.045 1.580 ;
        RECT 1.795 1.250 2.045 1.410 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.365 7.585 1.410 ;
        RECT 11.615 1.365 11.905 1.410 ;
        RECT 7.295 1.225 11.905 1.365 ;
        RECT 7.295 1.180 7.585 1.225 ;
        RECT 11.615 1.180 11.905 1.225 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 14.880 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.910 0.955 4.385 1.240 ;
        RECT 2.910 0.920 6.570 0.955 ;
        RECT 7.675 0.920 10.585 1.140 ;
        RECT 12.925 0.920 14.875 1.260 ;
        RECT 0.005 0.245 14.875 0.920 ;
        RECT 0.000 0.000 14.880 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 15.070 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 14.880 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 13.995 2.150 14.275 2.980 ;
        RECT 13.995 1.820 14.755 2.150 ;
        RECT 14.325 1.490 14.755 1.820 ;
        RECT 14.175 1.320 14.755 1.490 ;
        RECT 14.175 1.150 14.345 1.320 ;
        RECT 13.990 0.370 14.345 1.150 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 14.880 3.415 ;
        RECT 0.115 2.490 0.365 2.980 ;
        RECT 0.565 2.660 0.895 3.245 ;
        RECT 1.435 2.660 2.385 2.910 ;
        RECT 2.560 2.830 2.890 3.245 ;
        RECT 2.215 2.490 3.120 2.660 ;
        RECT 3.545 2.580 3.875 3.245 ;
        RECT 4.075 2.895 5.730 3.065 ;
        RECT 4.075 2.580 4.325 2.895 ;
        RECT 0.115 2.320 2.045 2.490 ;
        RECT 0.115 2.310 0.365 2.320 ;
        RECT 0.115 1.230 0.285 2.310 ;
        RECT 1.795 1.830 2.045 2.320 ;
        RECT 0.115 0.900 1.225 1.230 ;
        RECT 2.215 1.080 2.385 2.490 ;
        RECT 2.950 2.410 3.120 2.490 ;
        RECT 4.585 2.410 4.915 2.725 ;
        RECT 2.950 2.240 4.915 2.410 ;
        RECT 5.115 2.265 5.365 2.725 ;
        RECT 4.585 2.070 4.915 2.240 ;
        RECT 1.560 0.910 2.385 1.080 ;
        RECT 2.960 1.820 4.215 2.070 ;
        RECT 2.960 1.010 3.130 1.820 ;
        RECT 3.885 1.350 4.215 1.820 ;
        RECT 4.420 1.900 4.915 2.070 ;
        RECT 0.115 0.350 0.445 0.900 ;
        RECT 0.615 0.085 1.070 0.680 ;
        RECT 1.560 0.350 1.890 0.910 ;
        RECT 2.460 0.085 2.790 0.740 ;
        RECT 2.960 0.350 3.350 1.010 ;
        RECT 3.520 0.085 3.850 1.010 ;
        RECT 4.030 0.425 4.200 1.130 ;
        RECT 4.420 0.845 4.590 1.900 ;
        RECT 4.760 1.185 4.965 1.730 ;
        RECT 5.135 1.545 5.305 2.265 ;
        RECT 5.560 2.255 5.730 2.895 ;
        RECT 6.095 2.425 6.345 3.245 ;
        RECT 6.515 2.905 7.365 3.075 ;
        RECT 6.515 2.255 6.685 2.905 ;
        RECT 5.560 2.085 6.685 2.255 ;
        RECT 5.560 2.045 5.730 2.085 ;
        RECT 5.475 1.715 5.730 2.045 ;
        RECT 6.855 1.915 7.025 2.735 ;
        RECT 5.940 1.745 7.025 1.915 ;
        RECT 7.195 1.895 7.365 2.905 ;
        RECT 7.535 2.065 7.705 3.245 ;
        RECT 7.905 2.235 8.235 2.755 ;
        RECT 8.435 2.405 8.685 3.245 ;
        RECT 9.000 2.905 10.435 3.075 ;
        RECT 9.000 2.315 9.330 2.905 ;
        RECT 7.905 2.145 8.765 2.235 ;
        RECT 9.500 2.145 9.830 2.735 ;
        RECT 10.105 2.475 10.435 2.905 ;
        RECT 11.080 2.645 11.330 3.245 ;
        RECT 11.530 2.475 11.860 2.980 ;
        RECT 10.105 2.305 11.860 2.475 ;
        RECT 12.060 2.480 12.310 2.980 ;
        RECT 12.510 2.650 12.840 3.245 ;
        RECT 12.060 2.310 12.805 2.480 ;
        RECT 7.905 2.065 9.830 2.145 ;
        RECT 10.890 2.140 11.860 2.305 ;
        RECT 8.595 1.975 9.830 2.065 ;
        RECT 7.195 1.805 8.425 1.895 ;
        RECT 10.000 1.805 10.720 2.135 ;
        RECT 10.890 1.970 12.465 2.140 ;
        RECT 5.940 1.715 6.270 1.745 ;
        RECT 7.195 1.725 10.170 1.805 ;
        RECT 6.550 1.545 6.880 1.570 ;
        RECT 5.135 1.375 6.880 1.545 ;
        RECT 4.760 1.015 5.170 1.185 ;
        RECT 4.420 0.595 4.830 0.845 ;
        RECT 5.000 0.425 5.170 1.015 ;
        RECT 4.030 0.255 5.170 0.425 ;
        RECT 5.340 0.385 5.590 1.375 ;
        RECT 5.980 0.700 6.310 1.205 ;
        RECT 6.550 1.040 6.880 1.375 ;
        RECT 7.205 1.210 7.555 1.555 ;
        RECT 7.755 1.225 8.085 1.555 ;
        RECT 8.255 1.475 10.170 1.725 ;
        RECT 10.890 1.570 11.060 1.970 ;
        RECT 10.410 1.400 11.060 1.570 ;
        RECT 7.755 1.040 7.925 1.225 ;
        RECT 6.550 0.870 7.925 1.040 ;
        RECT 8.180 0.885 10.080 1.055 ;
        RECT 5.980 0.530 7.020 0.700 ;
        RECT 6.130 0.085 6.460 0.360 ;
        RECT 6.690 0.350 7.020 0.530 ;
        RECT 7.510 0.085 8.010 0.680 ;
        RECT 8.180 0.350 8.510 0.885 ;
        RECT 8.690 0.085 9.020 0.715 ;
        RECT 9.250 0.425 9.580 0.715 ;
        RECT 9.750 0.595 10.080 0.885 ;
        RECT 10.410 0.810 10.580 1.400 ;
        RECT 10.250 0.425 10.580 0.810 ;
        RECT 10.945 0.960 11.275 1.230 ;
        RECT 11.445 1.180 11.875 1.800 ;
        RECT 12.135 1.130 12.465 1.970 ;
        RECT 12.635 0.960 12.805 2.310 ;
        RECT 10.945 0.790 12.805 0.960 ;
        RECT 9.250 0.255 10.580 0.425 ;
        RECT 11.640 0.085 12.330 0.600 ;
        RECT 12.500 0.350 12.805 0.790 ;
        RECT 13.035 1.650 13.370 2.980 ;
        RECT 13.540 1.820 13.825 3.245 ;
        RECT 14.445 2.320 14.775 3.245 ;
        RECT 13.035 1.320 14.005 1.650 ;
        RECT 13.035 0.470 13.365 1.320 ;
        RECT 13.555 0.085 13.805 1.150 ;
        RECT 14.515 0.085 14.765 1.150 ;
        RECT 0.000 -0.085 14.880 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 7.355 1.210 7.525 1.380 ;
        RECT 11.675 1.210 11.845 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
  END
END sky130_fd_sc_hs__sdfstp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfstp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.345 1.180 3.715 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.105 1.820 1.575 2.150 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.100 2.835 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.580 0.855 2.150 ;
        RECT 0.525 1.410 2.045 1.580 ;
        RECT 1.715 1.250 2.045 1.410 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.735 7.585 1.780 ;
        RECT 11.615 1.735 11.905 1.780 ;
        RECT 7.295 1.595 11.905 1.735 ;
        RECT 7.295 1.550 7.585 1.595 ;
        RECT 11.615 1.550 11.905 1.595 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 15.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.950 1.035 4.430 1.240 ;
        RECT 12.770 1.210 15.730 1.240 ;
        RECT 2.950 0.955 4.990 1.035 ;
        RECT 2.950 0.920 6.650 0.955 ;
        RECT 7.725 0.920 10.650 1.140 ;
        RECT 12.770 0.920 15.835 1.210 ;
        RECT 0.005 0.245 15.835 0.920 ;
        RECT 0.000 0.000 15.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 15.840 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.201100 ;
    PORT
      LAYER li1 ;
        RECT 14.045 2.150 14.325 2.980 ;
        RECT 15.025 2.150 15.195 2.980 ;
        RECT 14.045 1.820 15.195 2.150 ;
        RECT 15.025 1.780 15.195 1.820 ;
        RECT 15.025 1.610 15.715 1.780 ;
        RECT 15.485 1.440 15.715 1.610 ;
        RECT 14.895 1.270 15.715 1.440 ;
        RECT 14.895 1.150 15.225 1.270 ;
        RECT 13.895 0.980 15.225 1.150 ;
        RECT 13.895 0.350 14.225 0.980 ;
        RECT 14.895 0.350 15.225 0.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 15.840 3.415 ;
        RECT 0.105 2.490 0.355 2.980 ;
        RECT 0.555 2.660 0.885 3.245 ;
        RECT 1.425 2.660 2.385 2.910 ;
        RECT 2.560 2.830 2.890 3.245 ;
        RECT 2.215 2.490 3.175 2.660 ;
        RECT 3.570 2.580 3.900 3.245 ;
        RECT 4.070 2.895 5.830 3.065 ;
        RECT 4.070 2.580 4.400 2.895 ;
        RECT 0.105 2.320 2.045 2.490 ;
        RECT 0.105 1.240 0.355 2.320 ;
        RECT 1.785 1.830 2.045 2.320 ;
        RECT 0.105 0.910 1.140 1.240 ;
        RECT 2.215 1.080 2.385 2.490 ;
        RECT 3.005 2.410 3.175 2.490 ;
        RECT 4.700 2.410 5.030 2.725 ;
        RECT 3.005 2.240 5.030 2.410 ;
        RECT 1.790 0.910 2.385 1.080 ;
        RECT 3.005 1.820 4.215 2.070 ;
        RECT 3.005 1.010 3.175 1.820 ;
        RECT 3.885 1.350 4.215 1.820 ;
        RECT 4.410 1.900 5.030 2.240 ;
        RECT 5.200 2.275 5.480 2.725 ;
        RECT 5.660 2.460 5.830 2.895 ;
        RECT 6.275 2.630 6.525 3.245 ;
        RECT 6.695 2.895 7.545 3.065 ;
        RECT 6.695 2.460 6.865 2.895 ;
        RECT 5.660 2.290 6.865 2.460 ;
        RECT 0.105 0.350 0.445 0.910 ;
        RECT 1.790 0.740 1.960 0.910 ;
        RECT 0.615 0.085 0.945 0.740 ;
        RECT 1.475 0.410 1.960 0.740 ;
        RECT 2.450 0.085 2.780 0.740 ;
        RECT 3.005 0.350 3.390 1.010 ;
        RECT 3.560 0.085 3.890 1.010 ;
        RECT 4.070 0.425 4.240 1.130 ;
        RECT 4.410 0.925 4.580 1.900 ;
        RECT 4.750 1.265 5.030 1.730 ;
        RECT 5.200 1.605 5.370 2.275 ;
        RECT 5.660 2.105 5.830 2.290 ;
        RECT 7.035 2.120 7.205 2.725 ;
        RECT 5.540 1.775 5.830 2.105 ;
        RECT 6.040 1.950 7.205 2.120 ;
        RECT 7.375 2.120 7.545 2.895 ;
        RECT 7.715 2.290 7.885 3.245 ;
        RECT 8.085 2.290 8.365 2.715 ;
        RECT 8.535 2.460 8.865 3.245 ;
        RECT 9.095 2.860 10.375 3.075 ;
        RECT 9.095 2.600 9.375 2.860 ;
        RECT 9.545 2.290 9.875 2.690 ;
        RECT 10.045 2.480 10.375 2.860 ;
        RECT 10.545 2.650 10.955 2.980 ;
        RECT 11.125 2.650 11.375 3.245 ;
        RECT 11.575 2.480 11.905 2.980 ;
        RECT 12.135 2.650 12.550 2.980 ;
        RECT 10.045 2.310 12.210 2.480 ;
        RECT 8.085 2.120 9.875 2.290 ;
        RECT 7.375 1.950 7.895 2.120 ;
        RECT 9.545 2.100 9.875 2.120 ;
        RECT 6.040 1.780 6.370 1.950 ;
        RECT 7.725 1.930 9.375 1.950 ;
        RECT 10.435 1.930 10.765 2.135 ;
        RECT 7.725 1.780 10.765 1.930 ;
        RECT 6.625 1.605 6.955 1.780 ;
        RECT 5.200 1.435 6.955 1.605 ;
        RECT 7.195 1.450 7.555 1.780 ;
        RECT 9.045 1.760 10.765 1.780 ;
        RECT 9.045 1.450 9.375 1.760 ;
        RECT 10.935 1.570 11.105 2.310 ;
        RECT 4.750 1.095 5.140 1.265 ;
        RECT 4.410 0.595 4.800 0.925 ;
        RECT 4.970 0.425 5.140 1.095 ;
        RECT 4.070 0.255 5.140 0.425 ;
        RECT 5.310 0.385 5.640 1.435 ;
        RECT 6.625 1.280 6.955 1.435 ;
        RECT 7.935 1.280 8.265 1.450 ;
        RECT 10.210 1.400 11.105 1.570 ;
        RECT 11.470 1.470 11.870 2.140 ;
        RECT 12.040 2.010 12.210 2.310 ;
        RECT 12.380 2.350 12.550 2.650 ;
        RECT 12.720 2.520 12.970 3.245 ;
        RECT 12.380 2.180 12.710 2.350 ;
        RECT 6.005 0.940 6.335 1.265 ;
        RECT 6.625 1.110 8.265 1.280 ;
        RECT 8.440 1.110 10.030 1.280 ;
        RECT 6.005 0.770 7.100 0.940 ;
        RECT 6.210 0.085 6.540 0.600 ;
        RECT 6.770 0.350 7.100 0.770 ;
        RECT 7.590 0.085 8.260 0.930 ;
        RECT 8.440 0.350 8.610 1.110 ;
        RECT 8.790 0.085 9.120 0.940 ;
        RECT 9.350 0.425 9.680 0.940 ;
        RECT 9.860 0.595 10.030 1.110 ;
        RECT 10.210 0.425 10.540 1.400 ;
        RECT 12.040 1.340 12.370 2.010 ;
        RECT 10.955 1.070 11.285 1.230 ;
        RECT 12.540 1.070 12.710 2.180 ;
        RECT 13.170 1.650 13.340 2.980 ;
        RECT 13.540 2.100 13.870 3.245 ;
        RECT 14.495 2.320 14.825 3.245 ;
        RECT 15.395 1.950 15.725 3.245 ;
        RECT 13.170 1.490 14.695 1.650 ;
        RECT 10.955 0.900 12.710 1.070 ;
        RECT 9.350 0.255 10.540 0.425 ;
        RECT 11.650 0.085 12.150 0.680 ;
        RECT 12.320 0.350 12.710 0.900 ;
        RECT 12.880 1.320 14.695 1.490 ;
        RECT 12.880 0.350 13.210 1.320 ;
        RECT 13.380 0.085 13.710 1.130 ;
        RECT 14.395 0.085 14.725 0.810 ;
        RECT 15.395 0.085 15.725 1.100 ;
        RECT 0.000 -0.085 15.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 7.355 1.580 7.525 1.750 ;
        RECT 11.675 1.580 11.845 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
  END
END sky130_fd_sc_hs__sdfstp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.235 1.180 3.685 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.455 1.630 1.785 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.380 1.550 2.725 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.955 2.050 1.285 ;
        RECT 1.565 0.810 2.050 0.955 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.480 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.530 1.050 4.540 1.240 ;
        RECT 9.960 1.050 12.475 1.240 ;
        RECT 2.530 0.920 8.025 1.050 ;
        RECT 8.970 0.920 12.475 1.050 ;
        RECT 0.025 0.245 12.475 0.920 ;
        RECT 0.000 0.000 12.480 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 12.670 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.480 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518900 ;
    PORT
      LAYER li1 ;
        RECT 10.650 1.820 10.915 2.980 ;
        RECT 10.745 1.130 10.915 1.820 ;
        RECT 10.500 0.350 10.915 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 12.045 1.820 12.375 2.980 ;
        RECT 12.155 1.050 12.375 1.820 ;
        RECT 12.035 0.350 12.375 1.050 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.480 3.415 ;
        RECT 0.085 1.855 0.530 2.980 ;
        RECT 0.700 2.300 1.030 3.245 ;
        RECT 1.570 2.560 1.900 2.980 ;
        RECT 2.560 2.730 3.150 3.245 ;
        RECT 3.830 2.730 4.335 3.245 ;
        RECT 4.985 2.630 5.235 2.920 ;
        RECT 4.505 2.560 5.235 2.630 ;
        RECT 1.570 2.460 5.235 2.560 ;
        RECT 5.410 2.460 5.765 2.920 ;
        RECT 6.450 2.860 6.780 3.245 ;
        RECT 5.935 2.520 7.735 2.690 ;
        RECT 1.570 2.390 4.675 2.460 ;
        RECT 1.570 2.300 1.900 2.390 ;
        RECT 0.745 1.955 2.170 2.125 ;
        RECT 0.745 1.855 0.915 1.955 ;
        RECT 0.085 1.525 0.915 1.855 ;
        RECT 1.840 1.795 2.170 1.955 ;
        RECT 0.085 0.785 0.255 1.525 ;
        RECT 2.895 1.350 3.065 2.390 ;
        RECT 3.270 1.990 3.600 2.220 ;
        RECT 3.270 1.820 4.025 1.990 ;
        RECT 2.220 1.180 3.065 1.350 ;
        RECT 0.085 0.350 0.465 0.785 ;
        RECT 0.635 0.085 0.965 0.730 ;
        RECT 2.220 0.640 2.390 1.180 ;
        RECT 3.855 1.010 4.025 1.820 ;
        RECT 4.195 1.650 4.365 2.390 ;
        RECT 4.910 2.220 5.240 2.280 ;
        RECT 4.535 1.820 5.240 2.220 ;
        RECT 4.195 1.480 4.900 1.650 ;
        RECT 3.035 0.840 4.025 1.010 ;
        RECT 1.455 0.390 2.390 0.640 ;
        RECT 2.615 0.085 2.865 0.810 ;
        RECT 3.035 0.350 3.365 0.840 ;
        RECT 3.595 0.085 3.935 0.670 ;
        RECT 4.195 0.425 4.445 1.130 ;
        RECT 4.650 0.595 4.900 1.480 ;
        RECT 5.070 0.425 5.240 1.820 ;
        RECT 5.410 1.700 5.580 2.460 ;
        RECT 5.935 2.200 6.105 2.520 ;
        RECT 5.750 1.870 6.105 2.200 ;
        RECT 6.985 2.100 7.395 2.350 ;
        RECT 6.690 1.700 7.020 1.930 ;
        RECT 5.410 1.530 7.020 1.700 ;
        RECT 5.410 0.595 5.580 1.530 ;
        RECT 7.190 1.360 7.360 2.100 ;
        RECT 7.565 1.960 7.735 2.520 ;
        RECT 7.905 2.130 8.235 2.980 ;
        RECT 8.860 2.650 9.430 3.245 ;
        RECT 9.600 2.350 9.950 2.980 ;
        RECT 7.565 1.630 7.880 1.960 ;
        RECT 8.065 1.950 8.235 2.130 ;
        RECT 8.710 2.120 9.950 2.350 ;
        RECT 8.065 1.780 9.020 1.950 ;
        RECT 9.600 1.940 9.950 2.120 ;
        RECT 8.050 1.420 8.680 1.610 ;
        RECT 5.750 0.860 6.035 1.360 ;
        RECT 6.245 1.030 7.360 1.360 ;
        RECT 7.530 1.355 8.680 1.420 ;
        RECT 7.530 1.250 8.220 1.355 ;
        RECT 8.850 1.270 9.020 1.780 ;
        RECT 9.280 1.270 9.610 1.770 ;
        RECT 7.530 1.090 7.860 1.250 ;
        RECT 8.850 1.150 9.610 1.270 ;
        RECT 7.190 0.920 7.360 1.030 ;
        RECT 5.750 0.690 7.020 0.860 ;
        RECT 5.750 0.425 6.035 0.690 ;
        RECT 4.195 0.255 6.035 0.425 ;
        RECT 6.430 0.085 6.680 0.520 ;
        RECT 6.850 0.425 7.020 0.690 ;
        RECT 7.190 0.595 7.520 0.920 ;
        RECT 7.690 0.425 7.860 1.090 ;
        RECT 8.390 1.100 9.610 1.150 ;
        RECT 9.780 1.650 9.950 1.940 ;
        RECT 10.120 1.820 10.450 3.245 ;
        RECT 9.780 1.320 10.575 1.650 ;
        RECT 11.090 1.550 11.340 2.875 ;
        RECT 11.540 1.995 11.870 3.245 ;
        RECT 8.390 0.980 9.020 1.100 ;
        RECT 8.390 0.810 8.560 0.980 ;
        RECT 9.780 0.930 9.950 1.320 ;
        RECT 11.090 1.220 11.985 1.550 ;
        RECT 6.850 0.255 7.860 0.425 ;
        RECT 8.030 0.350 8.560 0.810 ;
        RECT 8.740 0.085 9.410 0.810 ;
        RECT 9.590 0.350 9.950 0.930 ;
        RECT 10.150 0.085 10.320 1.130 ;
        RECT 11.090 0.540 11.310 1.220 ;
        RECT 11.490 0.085 11.865 1.020 ;
        RECT 0.000 -0.085 12.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
  END
END sky130_fd_sc_hs__sdfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.265 1.350 3.685 1.780 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.470 1.655 1.800 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.775 2.755 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.900 2.075 1.230 ;
        RECT 1.565 0.810 2.075 0.900 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 13.440 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 11.500 1.240 13.400 1.260 ;
        RECT 2.585 1.035 4.540 1.240 ;
        RECT 6.595 1.035 7.935 1.050 ;
        RECT 2.585 0.920 7.935 1.035 ;
        RECT 9.055 0.920 13.400 1.240 ;
        RECT 0.050 0.840 13.400 0.920 ;
        RECT 0.050 0.245 13.435 0.840 ;
        RECT 0.000 0.000 13.440 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 13.630 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 13.440 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 10.590 1.970 10.840 2.980 ;
        RECT 10.590 1.800 10.950 1.970 ;
        RECT 10.780 1.130 10.950 1.800 ;
        RECT 10.620 0.350 10.950 1.130 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.554300 ;
    PORT
      LAYER li1 ;
        RECT 12.555 2.150 12.835 2.980 ;
        RECT 12.555 1.820 13.315 2.150 ;
        RECT 13.075 1.150 13.315 1.820 ;
        RECT 12.550 0.900 13.315 1.150 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 13.440 3.415 ;
        RECT 0.085 1.800 0.520 2.925 ;
        RECT 0.725 2.310 1.055 3.245 ;
        RECT 1.650 2.540 1.980 2.925 ;
        RECT 2.670 2.710 3.090 3.245 ;
        RECT 4.075 2.710 4.405 3.245 ;
        RECT 6.575 2.955 6.905 3.245 ;
        RECT 5.085 2.665 5.335 2.935 ;
        RECT 4.575 2.540 5.335 2.665 ;
        RECT 1.650 2.495 5.335 2.540 ;
        RECT 1.650 2.370 4.745 2.495 ;
        RECT 5.505 2.475 5.865 2.935 ;
        RECT 6.035 2.615 7.735 2.785 ;
        RECT 1.650 2.310 1.980 2.370 ;
        RECT 0.745 1.970 2.195 2.140 ;
        RECT 0.745 1.800 0.915 1.970 ;
        RECT 0.085 1.470 0.915 1.800 ;
        RECT 1.865 1.725 2.195 1.970 ;
        RECT 2.925 1.520 3.095 2.370 ;
        RECT 3.295 1.950 4.095 2.200 ;
        RECT 0.085 0.730 0.255 1.470 ;
        RECT 2.245 1.350 3.095 1.520 ;
        RECT 3.855 1.350 4.095 1.950 ;
        RECT 4.265 1.650 4.435 2.370 ;
        RECT 5.005 2.200 5.335 2.325 ;
        RECT 4.605 2.005 5.335 2.200 ;
        RECT 4.605 1.820 4.855 2.005 ;
        RECT 4.265 1.480 4.900 1.650 ;
        RECT 0.085 0.350 0.490 0.730 ;
        RECT 0.660 0.085 0.990 0.730 ;
        RECT 2.245 0.640 2.415 1.350 ;
        RECT 3.855 1.180 4.025 1.350 ;
        RECT 1.480 0.390 2.415 0.640 ;
        RECT 2.695 0.085 2.945 1.130 ;
        RECT 3.125 1.010 4.025 1.180 ;
        RECT 3.125 0.350 3.455 1.010 ;
        RECT 3.685 0.085 4.015 0.840 ;
        RECT 4.195 0.425 4.445 1.130 ;
        RECT 4.650 0.595 4.900 1.480 ;
        RECT 5.070 0.425 5.240 2.005 ;
        RECT 5.505 1.745 5.675 2.475 ;
        RECT 6.035 2.245 6.205 2.615 ;
        RECT 5.845 1.915 6.205 2.245 ;
        RECT 7.110 2.115 7.395 2.445 ;
        RECT 6.730 1.745 7.010 1.945 ;
        RECT 5.410 1.575 7.010 1.745 ;
        RECT 5.410 0.875 5.580 1.575 ;
        RECT 7.180 1.405 7.350 2.115 ;
        RECT 7.565 1.930 7.735 2.615 ;
        RECT 7.905 2.100 8.235 2.980 ;
        RECT 8.860 2.650 9.430 3.245 ;
        RECT 9.600 2.380 9.950 2.980 ;
        RECT 7.565 1.600 7.895 1.930 ;
        RECT 8.065 1.890 8.235 2.100 ;
        RECT 8.710 2.060 9.950 2.380 ;
        RECT 9.600 1.940 9.950 2.060 ;
        RECT 8.065 1.720 9.020 1.890 ;
        RECT 5.750 1.045 6.080 1.375 ;
        RECT 6.250 1.110 7.350 1.405 ;
        RECT 8.350 1.395 8.680 1.550 ;
        RECT 5.910 0.940 6.080 1.045 ;
        RECT 5.410 0.595 5.740 0.875 ;
        RECT 5.910 0.770 7.010 0.940 ;
        RECT 5.910 0.425 6.080 0.770 ;
        RECT 4.195 0.255 6.080 0.425 ;
        RECT 6.340 0.085 6.670 0.600 ;
        RECT 6.840 0.425 7.010 0.770 ;
        RECT 7.180 0.595 7.350 1.110 ;
        RECT 7.520 1.225 8.680 1.395 ;
        RECT 8.850 1.225 9.020 1.720 ;
        RECT 9.780 1.630 9.950 1.940 ;
        RECT 10.140 1.820 10.390 3.245 ;
        RECT 11.040 2.140 11.370 3.245 ;
        RECT 11.120 1.820 11.370 2.140 ;
        RECT 11.580 1.650 11.910 2.860 ;
        RECT 12.105 1.820 12.355 3.245 ;
        RECT 13.005 2.320 13.335 3.245 ;
        RECT 9.280 1.225 9.610 1.550 ;
        RECT 7.520 1.030 7.780 1.225 ;
        RECT 8.850 1.055 9.610 1.225 ;
        RECT 9.780 1.300 10.610 1.630 ;
        RECT 11.580 1.320 12.735 1.650 ;
        RECT 7.520 0.425 7.690 1.030 ;
        RECT 8.020 0.885 9.020 1.055 ;
        RECT 9.780 0.885 9.950 1.300 ;
        RECT 8.020 0.810 8.190 0.885 ;
        RECT 6.840 0.255 7.690 0.425 ;
        RECT 7.860 0.350 8.190 0.810 ;
        RECT 8.680 0.085 9.390 0.715 ;
        RECT 9.560 0.350 9.950 0.885 ;
        RECT 10.120 0.085 10.450 1.130 ;
        RECT 11.130 0.085 11.380 1.130 ;
        RECT 11.580 0.560 11.940 1.320 ;
        RECT 12.120 0.730 12.380 1.150 ;
        RECT 12.120 0.085 12.450 0.730 ;
        RECT 12.995 0.085 13.325 0.730 ;
        RECT 0.000 -0.085 13.440 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
  END
END sky130_fd_sc_hs__sdfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.250 1.180 3.685 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.455 1.655 1.785 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.470 2.740 2.140 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.955 2.250 1.285 ;
        RECT 1.085 0.900 2.250 0.955 ;
        RECT 1.085 0.810 1.315 0.900 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 11.040 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.585 1.050 4.535 1.240 ;
        RECT 10.080 1.050 11.035 1.260 ;
        RECT 2.585 0.920 11.035 1.050 ;
        RECT 0.045 0.245 11.035 0.920 ;
        RECT 0.000 0.000 11.040 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 11.230 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 11.040 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.528300 ;
    PORT
      LAYER li1 ;
        RECT 10.600 0.370 10.935 2.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 11.040 3.415 ;
        RECT 0.085 2.125 0.555 2.980 ;
        RECT 0.725 2.300 1.055 3.245 ;
        RECT 1.595 2.480 1.925 2.980 ;
        RECT 2.670 2.650 3.175 3.245 ;
        RECT 3.855 2.730 4.365 3.245 ;
        RECT 4.535 2.710 5.375 2.980 ;
        RECT 4.535 2.560 4.705 2.710 ;
        RECT 3.345 2.480 4.705 2.560 ;
        RECT 5.545 2.540 5.875 2.980 ;
        RECT 6.480 2.860 6.810 3.245 ;
        RECT 1.595 2.390 4.705 2.480 ;
        RECT 1.595 2.310 4.395 2.390 ;
        RECT 1.865 2.125 2.195 2.140 ;
        RECT 0.085 1.955 2.195 2.125 ;
        RECT 0.085 1.525 0.825 1.955 ;
        RECT 0.085 0.785 0.255 1.525 ;
        RECT 1.865 1.470 2.195 1.955 ;
        RECT 2.910 1.300 3.080 2.310 ;
        RECT 3.295 1.820 4.055 2.140 ;
        RECT 2.420 1.130 3.080 1.300 ;
        RECT 3.855 1.300 4.055 1.820 ;
        RECT 4.225 1.650 4.395 2.310 ;
        RECT 4.955 2.220 5.225 2.380 ;
        RECT 4.565 2.050 5.225 2.220 ;
        RECT 4.565 1.820 4.815 2.050 ;
        RECT 4.225 1.480 4.785 1.650 ;
        RECT 0.085 0.350 0.405 0.785 ;
        RECT 0.585 0.085 0.915 0.785 ;
        RECT 2.420 0.730 2.590 1.130 ;
        RECT 3.855 0.960 4.025 1.300 ;
        RECT 3.125 0.790 4.025 0.960 ;
        RECT 1.485 0.400 2.590 0.730 ;
        RECT 2.775 0.085 2.945 0.790 ;
        RECT 3.125 0.350 3.455 0.790 ;
        RECT 3.685 0.085 4.015 0.620 ;
        RECT 4.195 0.425 4.445 1.130 ;
        RECT 4.615 0.940 4.785 1.480 ;
        RECT 4.615 0.595 4.885 0.940 ;
        RECT 5.055 0.425 5.225 2.050 ;
        RECT 5.395 2.370 5.875 2.540 ;
        RECT 6.045 2.520 7.715 2.690 ;
        RECT 5.395 1.700 5.565 2.370 ;
        RECT 6.045 2.200 6.215 2.520 ;
        RECT 5.735 1.870 6.215 2.200 ;
        RECT 7.015 2.100 7.375 2.350 ;
        RECT 6.645 1.700 6.975 1.930 ;
        RECT 5.395 1.530 6.975 1.700 ;
        RECT 5.395 0.595 5.565 1.530 ;
        RECT 7.145 1.360 7.315 2.100 ;
        RECT 7.545 1.930 7.715 2.520 ;
        RECT 7.885 2.415 8.135 2.980 ;
        RECT 8.845 2.650 9.420 3.245 ;
        RECT 7.885 2.245 8.895 2.415 ;
        RECT 7.885 2.100 8.135 2.245 ;
        RECT 7.545 1.600 7.900 1.930 ;
        RECT 8.305 1.490 8.555 2.075 ;
        RECT 8.070 1.360 8.555 1.490 ;
        RECT 5.735 0.860 5.985 1.360 ;
        RECT 6.195 1.030 7.315 1.360 ;
        RECT 7.485 1.320 8.555 1.360 ;
        RECT 8.725 1.930 8.895 2.245 ;
        RECT 9.590 2.100 9.935 2.980 ;
        RECT 8.725 1.600 9.595 1.930 ;
        RECT 9.765 1.650 9.935 2.100 ;
        RECT 10.150 1.820 10.400 3.245 ;
        RECT 7.485 1.190 8.240 1.320 ;
        RECT 7.485 1.030 7.815 1.190 ;
        RECT 8.725 1.150 8.895 1.600 ;
        RECT 9.765 1.360 10.245 1.650 ;
        RECT 7.145 0.860 7.315 1.030 ;
        RECT 5.735 0.690 6.975 0.860 ;
        RECT 5.735 0.425 5.905 0.690 ;
        RECT 4.195 0.255 5.905 0.425 ;
        RECT 6.385 0.085 6.635 0.520 ;
        RECT 6.805 0.425 6.975 0.690 ;
        RECT 7.145 0.595 7.475 0.860 ;
        RECT 7.645 0.425 7.815 1.030 ;
        RECT 8.410 0.980 8.895 1.150 ;
        RECT 9.065 1.320 10.245 1.360 ;
        RECT 9.065 1.030 9.980 1.320 ;
        RECT 8.410 0.940 8.580 0.980 ;
        RECT 7.985 0.770 8.580 0.940 ;
        RECT 7.985 0.480 8.315 0.770 ;
        RECT 6.805 0.255 7.815 0.425 ;
        RECT 8.805 0.085 9.480 0.810 ;
        RECT 9.650 0.350 9.980 1.030 ;
        RECT 10.175 0.085 10.425 1.150 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
  END
END sky130_fd_sc_hs__sdfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.290 1.350 3.685 1.780 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.190 1.665 1.845 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.450 1.435 2.780 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.020 0.835 1.230 ;
        RECT 1.875 1.020 2.205 1.230 ;
        RECT 0.425 0.850 2.205 1.020 ;
        RECT 0.425 0.810 0.835 0.850 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.000 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.605 1.050 4.645 1.240 ;
        RECT 9.295 1.050 11.995 1.240 ;
        RECT 2.605 0.920 11.995 1.050 ;
        RECT 0.005 0.245 11.995 0.920 ;
        RECT 0.000 0.000 12.000 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 12.190 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.000 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.576500 ;
    PORT
      LAYER li1 ;
        RECT 11.105 1.820 11.435 2.980 ;
        RECT 11.215 1.050 11.385 1.820 ;
        RECT 11.055 0.350 11.385 1.050 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.000 3.415 ;
        RECT 0.085 2.185 0.445 2.925 ;
        RECT 0.615 2.355 0.945 3.245 ;
        RECT 1.485 2.620 2.060 2.945 ;
        RECT 2.685 2.790 3.135 3.245 ;
        RECT 3.900 2.790 4.370 3.245 ;
        RECT 5.135 2.620 5.385 2.980 ;
        RECT 1.485 2.450 5.385 2.620 ;
        RECT 5.555 2.520 5.915 2.980 ;
        RECT 6.585 2.520 6.835 3.245 ;
        RECT 7.005 2.905 7.855 3.075 ;
        RECT 1.485 2.355 3.120 2.450 ;
        RECT 0.085 2.015 2.210 2.185 ;
        RECT 0.085 1.470 0.915 2.015 ;
        RECT 1.880 1.775 2.210 2.015 ;
        RECT 0.085 0.640 0.255 1.470 ;
        RECT 2.950 1.265 3.120 2.355 ;
        RECT 3.340 1.950 4.145 2.280 ;
        RECT 2.375 1.095 3.120 1.265 ;
        RECT 3.855 1.300 4.145 1.950 ;
        RECT 4.315 1.470 4.485 2.450 ;
        RECT 4.655 1.820 5.375 2.280 ;
        RECT 5.045 1.610 5.375 1.820 ;
        RECT 5.555 1.800 5.725 2.520 ;
        RECT 7.005 2.300 7.175 2.905 ;
        RECT 5.895 2.130 7.175 2.300 ;
        RECT 5.895 1.970 6.225 2.130 ;
        RECT 6.845 1.800 7.175 1.960 ;
        RECT 5.555 1.630 7.175 1.800 ;
        RECT 4.315 1.300 4.875 1.470 ;
        RECT 3.855 1.180 4.025 1.300 ;
        RECT 2.375 0.680 2.545 1.095 ;
        RECT 3.305 1.010 4.025 1.180 ;
        RECT 3.305 0.920 3.475 1.010 ;
        RECT 0.085 0.390 0.490 0.640 ;
        RECT 0.660 0.085 0.990 0.640 ;
        RECT 1.480 0.350 2.545 0.680 ;
        RECT 2.715 0.085 2.975 0.810 ;
        RECT 3.145 0.330 3.475 0.920 ;
        RECT 3.705 0.085 4.035 0.840 ;
        RECT 4.205 0.425 4.535 1.130 ;
        RECT 4.705 0.940 4.875 1.300 ;
        RECT 4.705 0.595 5.015 0.940 ;
        RECT 5.185 0.425 5.355 1.610 ;
        RECT 5.555 0.940 5.775 1.630 ;
        RECT 7.345 1.390 7.515 2.610 ;
        RECT 7.685 1.930 7.855 2.905 ;
        RECT 8.025 2.660 8.275 2.920 ;
        RECT 8.025 2.490 9.060 2.660 ;
        RECT 9.295 2.590 9.925 3.245 ;
        RECT 8.285 1.990 8.720 2.320 ;
        RECT 8.890 2.245 9.060 2.490 ;
        RECT 10.095 2.415 10.445 2.920 ;
        RECT 8.890 2.075 10.105 2.245 ;
        RECT 7.685 1.600 8.115 1.930 ;
        RECT 5.525 0.595 5.775 0.940 ;
        RECT 5.945 0.890 6.275 1.360 ;
        RECT 6.485 1.230 7.515 1.390 ;
        RECT 8.285 1.360 8.455 1.990 ;
        RECT 6.485 1.060 7.890 1.230 ;
        RECT 5.945 0.720 7.390 0.890 ;
        RECT 5.945 0.425 6.115 0.720 ;
        RECT 4.205 0.255 6.115 0.425 ;
        RECT 6.720 0.085 7.050 0.550 ;
        RECT 7.220 0.425 7.390 0.720 ;
        RECT 7.560 0.595 7.890 1.060 ;
        RECT 8.060 1.030 8.455 1.360 ;
        RECT 8.060 0.425 8.230 1.030 ;
        RECT 8.890 0.810 9.060 2.075 ;
        RECT 9.230 1.240 9.535 1.905 ;
        RECT 9.775 1.410 10.105 2.075 ;
        RECT 10.275 1.550 10.445 2.415 ;
        RECT 10.655 1.820 10.905 3.245 ;
        RECT 11.635 1.820 11.885 3.245 ;
        RECT 10.275 1.240 11.045 1.550 ;
        RECT 9.230 1.220 11.045 1.240 ;
        RECT 9.230 1.070 10.445 1.220 ;
        RECT 7.220 0.255 8.230 0.425 ;
        RECT 8.400 0.640 9.060 0.810 ;
        RECT 8.400 0.350 8.795 0.640 ;
        RECT 9.300 0.085 9.630 0.810 ;
        RECT 9.800 0.350 10.130 1.070 ;
        RECT 10.615 0.085 10.885 1.050 ;
        RECT 11.555 0.085 11.885 1.130 ;
        RECT 0.000 -0.085 12.000 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
  END
END sky130_fd_sc_hs__sdfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 3.275 1.180 3.685 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.455 1.655 1.785 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.550 2.765 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.955 2.195 1.285 ;
        RECT 1.565 0.810 2.195 0.955 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 12.480 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.620 1.050 4.555 1.240 ;
        RECT 2.620 0.920 8.735 1.050 ;
        RECT 9.645 0.920 12.475 1.240 ;
        RECT 0.050 0.245 12.475 0.920 ;
        RECT 0.000 0.000 12.480 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 12.670 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 12.480 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.149300 ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.970 11.015 2.980 ;
        RECT 11.665 2.015 11.855 2.980 ;
        RECT 11.665 1.970 12.355 2.015 ;
        RECT 10.685 1.800 12.355 1.970 ;
        RECT 11.760 1.130 12.355 1.800 ;
        RECT 10.745 0.880 12.355 1.130 ;
        RECT 10.745 0.350 10.995 0.880 ;
        RECT 11.675 0.350 11.865 0.880 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 12.480 3.415 ;
        RECT 0.085 2.125 0.555 2.980 ;
        RECT 0.725 2.300 1.055 3.245 ;
        RECT 1.595 2.560 1.925 2.980 ;
        RECT 2.585 2.730 3.205 3.245 ;
        RECT 3.885 2.730 4.475 3.245 ;
        RECT 5.155 2.710 5.405 2.970 ;
        RECT 4.645 2.560 5.405 2.710 ;
        RECT 1.595 2.540 5.405 2.560 ;
        RECT 1.595 2.390 4.815 2.540 ;
        RECT 5.575 2.510 5.935 2.970 ;
        RECT 6.680 2.855 7.010 3.245 ;
        RECT 6.105 2.515 8.100 2.685 ;
        RECT 1.595 2.310 1.925 2.390 ;
        RECT 1.865 2.125 2.195 2.140 ;
        RECT 0.085 1.955 2.195 2.125 ;
        RECT 0.085 1.525 0.915 1.955 ;
        RECT 0.085 0.785 0.255 1.525 ;
        RECT 1.865 1.470 2.195 1.955 ;
        RECT 2.935 1.350 3.105 2.390 ;
        RECT 3.325 1.990 3.655 2.220 ;
        RECT 3.325 1.820 4.165 1.990 ;
        RECT 2.365 1.180 3.105 1.350 ;
        RECT 3.855 1.300 4.165 1.820 ;
        RECT 4.335 1.650 4.505 2.390 ;
        RECT 5.075 2.220 5.405 2.370 ;
        RECT 4.675 2.040 5.405 2.220 ;
        RECT 4.675 1.820 4.925 2.040 ;
        RECT 4.335 1.480 4.925 1.650 ;
        RECT 0.085 0.350 0.490 0.785 ;
        RECT 0.660 0.085 0.990 0.785 ;
        RECT 2.365 0.640 2.535 1.180 ;
        RECT 3.855 1.010 4.025 1.300 ;
        RECT 3.125 0.840 4.025 1.010 ;
        RECT 1.480 0.390 2.535 0.640 ;
        RECT 2.705 0.085 2.955 0.810 ;
        RECT 3.125 0.350 3.455 0.840 ;
        RECT 3.685 0.085 4.015 0.670 ;
        RECT 4.195 0.425 4.445 1.130 ;
        RECT 4.675 0.595 4.925 1.480 ;
        RECT 5.095 0.425 5.265 2.040 ;
        RECT 5.575 1.780 5.745 2.510 ;
        RECT 6.105 2.280 6.275 2.515 ;
        RECT 5.915 1.950 6.275 2.280 ;
        RECT 7.215 2.175 7.760 2.345 ;
        RECT 6.835 1.780 7.160 1.940 ;
        RECT 5.435 1.610 7.160 1.780 ;
        RECT 5.435 0.595 5.605 1.610 ;
        RECT 7.330 1.440 7.500 2.175 ;
        RECT 7.930 1.955 8.100 2.515 ;
        RECT 8.270 2.190 8.600 2.820 ;
        RECT 9.225 2.360 9.555 3.245 ;
        RECT 8.270 2.020 9.185 2.190 ;
        RECT 7.770 1.625 8.100 1.955 ;
        RECT 9.015 1.800 9.185 2.020 ;
        RECT 9.730 1.970 10.135 2.820 ;
        RECT 5.775 0.940 6.075 1.360 ;
        RECT 6.295 1.110 7.500 1.440 ;
        RECT 8.535 1.410 8.845 1.715 ;
        RECT 5.775 0.770 7.160 0.940 ;
        RECT 5.775 0.425 5.945 0.770 ;
        RECT 4.195 0.255 5.945 0.425 ;
        RECT 6.490 0.085 6.820 0.600 ;
        RECT 6.990 0.465 7.160 0.770 ;
        RECT 7.330 0.885 7.500 1.110 ;
        RECT 7.670 1.240 8.845 1.410 ;
        RECT 9.015 1.470 9.795 1.800 ;
        RECT 9.965 1.630 10.135 1.970 ;
        RECT 10.305 1.940 10.475 3.245 ;
        RECT 11.215 2.140 11.465 3.245 ;
        RECT 12.035 2.185 12.365 3.245 ;
        RECT 7.670 1.055 8.125 1.240 ;
        RECT 9.015 1.070 9.185 1.470 ;
        RECT 9.965 1.300 11.545 1.630 ;
        RECT 7.330 0.635 7.785 0.885 ;
        RECT 7.955 0.465 8.125 1.055 ;
        RECT 6.990 0.295 8.125 0.465 ;
        RECT 8.295 0.900 9.185 1.070 ;
        RECT 9.355 1.130 10.135 1.300 ;
        RECT 9.355 0.900 9.665 1.130 ;
        RECT 8.295 0.350 8.625 0.900 ;
        RECT 9.195 0.085 9.525 0.730 ;
        RECT 9.835 0.350 10.005 1.130 ;
        RECT 10.185 0.085 10.515 0.960 ;
        RECT 11.175 0.085 11.505 0.710 ;
        RECT 12.035 0.085 12.365 0.710 ;
        RECT 0.000 -0.085 12.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
  END
END sky130_fd_sc_hs__sdfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.680 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.459000 ;
    PORT
      LAYER li1 ;
        RECT 5.330 1.355 5.660 1.780 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.630 1.285 2.150 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.290 0.545 1.960 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 7.680 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.050 2.005 1.240 ;
        RECT 3.845 1.050 7.675 1.240 ;
        RECT 0.005 0.245 7.675 1.050 ;
        RECT 0.000 0.000 7.680 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 7.870 3.520 ;
        RECT 3.910 1.580 4.980 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 7.680 3.575 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632800 ;
    PORT
      LAYER li1 ;
        RECT 7.235 1.820 7.585 2.980 ;
        RECT 7.415 1.130 7.585 1.820 ;
        RECT 7.240 0.350 7.585 1.130 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 7.680 3.415 ;
        RECT 0.115 2.130 0.445 3.245 ;
        RECT 0.955 2.490 1.285 2.980 ;
        RECT 1.515 2.660 1.845 3.245 ;
        RECT 2.610 2.490 2.860 2.755 ;
        RECT 0.955 2.320 2.860 2.490 ;
        RECT 3.060 2.425 3.390 2.755 ;
        RECT 3.985 2.440 4.315 3.245 ;
        RECT 4.490 2.665 4.820 2.900 ;
        RECT 5.585 2.835 5.990 3.245 ;
        RECT 4.490 2.495 6.000 2.665 ;
        RECT 1.455 1.460 1.625 2.320 ;
        RECT 0.715 1.290 1.625 1.460 ;
        RECT 1.795 1.715 2.380 2.150 ;
        RECT 2.610 1.885 2.860 2.320 ;
        RECT 1.795 1.545 2.900 1.715 ;
        RECT 0.715 1.120 0.885 1.290 ;
        RECT 1.795 1.120 1.965 1.545 ;
        RECT 2.625 1.385 2.900 1.545 ;
        RECT 3.070 1.550 3.390 2.425 ;
        RECT 4.490 2.120 4.820 2.495 ;
        RECT 3.600 1.740 4.820 2.120 ;
        RECT 4.990 1.995 5.380 2.325 ;
        RECT 0.115 0.085 0.365 1.120 ;
        RECT 0.545 0.710 0.885 1.120 ;
        RECT 1.565 0.950 1.965 1.120 ;
        RECT 2.135 1.200 2.415 1.360 ;
        RECT 3.070 1.220 4.320 1.550 ;
        RECT 2.135 1.030 2.715 1.200 ;
        RECT 1.565 0.880 1.895 0.950 ;
        RECT 2.125 0.710 2.375 0.780 ;
        RECT 0.545 0.540 2.375 0.710 ;
        RECT 1.055 0.085 1.385 0.370 ;
        RECT 2.125 0.350 2.375 0.540 ;
        RECT 2.545 0.425 2.715 1.030 ;
        RECT 3.070 0.925 3.240 1.220 ;
        RECT 4.490 1.050 4.680 1.740 ;
        RECT 4.990 1.130 5.160 1.995 ;
        RECT 5.830 1.550 6.000 2.495 ;
        RECT 6.195 1.890 6.525 2.875 ;
        RECT 6.695 2.060 7.025 3.245 ;
        RECT 6.195 1.720 6.645 1.890 ;
        RECT 6.475 1.630 6.645 1.720 ;
        RECT 5.830 1.220 6.305 1.550 ;
        RECT 6.475 1.300 7.245 1.630 ;
        RECT 2.885 0.595 3.240 0.925 ;
        RECT 3.410 0.880 4.260 1.050 ;
        RECT 3.410 0.425 3.580 0.880 ;
        RECT 2.545 0.255 3.580 0.425 ;
        RECT 3.750 0.085 3.920 0.710 ;
        RECT 4.090 0.425 4.260 0.880 ;
        RECT 4.430 0.595 4.680 1.050 ;
        RECT 4.900 0.425 5.230 1.130 ;
        RECT 4.090 0.255 5.230 0.425 ;
        RECT 5.410 0.085 5.660 1.130 ;
        RECT 6.475 1.050 6.645 1.300 ;
        RECT 6.165 0.450 6.645 1.050 ;
        RECT 6.815 0.085 7.065 1.130 ;
        RECT 0.000 -0.085 7.680 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
  END
END sky130_fd_sc_hs__sdlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdlclkp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.498000 ;
    PORT
      LAYER li1 ;
        RECT 5.335 1.180 5.665 1.550 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.795 1.630 1.300 2.150 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.290 0.550 1.960 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.965 1.240 4.910 1.275 ;
        RECT 0.005 1.050 2.005 1.240 ;
        RECT 3.965 1.050 8.155 1.240 ;
        RECT 0.005 0.245 8.155 1.050 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
        RECT 3.840 1.560 5.890 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 7.210 1.820 7.565 2.980 ;
        RECT 7.395 1.130 7.565 1.820 ;
        RECT 7.295 0.350 7.625 1.130 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.105 2.130 0.435 3.245 ;
        RECT 0.945 2.490 1.275 2.980 ;
        RECT 1.485 2.660 1.815 3.245 ;
        RECT 2.550 2.490 2.800 2.755 ;
        RECT 0.945 2.320 2.800 2.490 ;
        RECT 1.470 1.390 1.640 2.320 ;
        RECT 0.720 1.220 1.640 1.390 ;
        RECT 1.810 1.715 2.340 2.150 ;
        RECT 2.550 1.885 2.800 2.320 ;
        RECT 3.000 2.235 3.360 2.695 ;
        RECT 1.810 1.545 3.020 1.715 ;
        RECT 0.720 1.120 0.890 1.220 ;
        RECT 0.115 0.085 0.365 1.120 ;
        RECT 0.545 0.710 0.890 1.120 ;
        RECT 1.810 1.050 1.980 1.545 ;
        RECT 2.690 1.385 3.020 1.545 ;
        RECT 3.190 1.415 3.360 2.235 ;
        RECT 3.990 2.095 4.240 3.245 ;
        RECT 4.440 2.390 4.825 2.920 ;
        RECT 5.510 2.560 5.840 3.245 ;
        RECT 4.440 2.220 6.005 2.390 ;
        RECT 4.440 1.925 4.825 2.220 ;
        RECT 3.530 1.755 4.825 1.925 ;
        RECT 3.530 1.585 3.860 1.755 ;
        RECT 4.155 1.415 4.485 1.585 ;
        RECT 1.565 0.880 1.980 1.050 ;
        RECT 2.150 1.200 2.480 1.360 ;
        RECT 3.190 1.245 4.485 1.415 ;
        RECT 2.150 1.030 2.715 1.200 ;
        RECT 0.545 0.540 2.375 0.710 ;
        RECT 1.055 0.085 1.385 0.370 ;
        RECT 2.125 0.350 2.375 0.540 ;
        RECT 2.545 0.425 2.715 1.030 ;
        RECT 3.190 0.845 3.360 1.245 ;
        RECT 4.655 1.075 4.825 1.755 ;
        RECT 2.885 0.595 3.360 0.845 ;
        RECT 3.530 0.905 4.380 1.075 ;
        RECT 3.530 0.425 3.700 0.905 ;
        RECT 2.545 0.255 3.700 0.425 ;
        RECT 3.870 0.085 4.040 0.735 ;
        RECT 4.210 0.425 4.380 0.905 ;
        RECT 4.550 0.595 4.825 1.075 ;
        RECT 4.995 1.720 5.310 2.050 ;
        RECT 4.995 1.010 5.165 1.720 ;
        RECT 5.835 1.630 6.005 2.220 ;
        RECT 6.175 1.970 6.505 2.890 ;
        RECT 6.710 2.140 7.040 3.245 ;
        RECT 6.175 1.800 7.040 1.970 ;
        RECT 7.740 1.820 7.990 3.245 ;
        RECT 6.870 1.630 7.040 1.800 ;
        RECT 5.835 1.300 6.530 1.630 ;
        RECT 6.870 1.300 7.225 1.630 ;
        RECT 6.870 1.130 7.040 1.300 ;
        RECT 4.995 0.425 5.360 1.010 ;
        RECT 4.210 0.255 5.360 0.425 ;
        RECT 5.530 0.085 5.860 1.010 ;
        RECT 6.325 0.960 7.040 1.130 ;
        RECT 6.325 0.350 6.655 0.960 ;
        RECT 6.865 0.085 7.115 0.790 ;
        RECT 7.805 0.085 8.055 1.130 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
  END
END sky130_fd_sc_hs__sdlclkp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdlclkp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.516000 ;
    PORT
      LAYER li1 ;
        RECT 5.785 1.180 6.115 1.550 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.455 1.315 1.785 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.208500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.455 0.550 1.785 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.050 2.185 1.395 ;
        RECT 4.440 1.050 9.595 1.240 ;
        RECT 0.005 0.245 9.595 1.050 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
        RECT 1.385 1.650 5.370 1.660 ;
        RECT 4.270 1.575 5.370 1.650 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.319400 ;
    PORT
      LAYER li1 ;
        RECT 7.705 1.970 8.035 2.980 ;
        RECT 8.655 1.970 8.985 2.980 ;
        RECT 7.705 1.800 8.985 1.970 ;
        RECT 8.725 1.410 8.985 1.800 ;
        RECT 8.725 1.130 9.055 1.410 ;
        RECT 7.865 0.960 9.055 1.130 ;
        RECT 7.865 0.350 8.115 0.960 ;
        RECT 8.725 0.350 9.055 0.960 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.115 1.955 0.445 3.245 ;
        RECT 0.985 2.480 1.315 2.835 ;
        RECT 1.545 2.650 2.160 3.245 ;
        RECT 2.925 2.480 3.255 2.755 ;
        RECT 0.985 2.310 3.255 2.480 ;
        RECT 0.985 1.955 1.655 2.310 ;
        RECT 0.115 0.085 0.445 1.285 ;
        RECT 0.615 0.785 0.945 1.285 ;
        RECT 1.485 0.785 1.655 1.955 ;
        RECT 2.365 1.735 2.695 2.140 ;
        RECT 2.925 1.905 3.255 2.310 ;
        RECT 1.825 1.565 3.255 1.735 ;
        RECT 1.825 0.955 2.075 1.565 ;
        RECT 2.925 1.405 3.255 1.565 ;
        RECT 3.425 1.405 3.705 2.755 ;
        RECT 4.430 2.075 4.680 3.245 ;
        RECT 4.880 2.410 5.270 2.895 ;
        RECT 5.980 2.580 6.310 3.245 ;
        RECT 4.880 2.240 6.455 2.410 ;
        RECT 4.880 1.905 5.270 2.240 ;
        RECT 3.960 1.735 5.270 1.905 ;
        RECT 5.440 1.820 5.775 2.070 ;
        RECT 3.960 1.575 4.290 1.735 ;
        RECT 4.600 1.405 4.930 1.565 ;
        RECT 2.245 1.235 2.575 1.395 ;
        RECT 3.425 1.235 4.930 1.405 ;
        RECT 2.245 1.065 2.975 1.235 ;
        RECT 2.305 0.785 2.635 0.895 ;
        RECT 0.615 0.615 2.635 0.785 ;
        RECT 1.125 0.085 1.565 0.445 ;
        RECT 2.305 0.350 2.635 0.615 ;
        RECT 2.805 0.440 2.975 1.065 ;
        RECT 3.425 0.940 3.595 1.235 ;
        RECT 5.100 1.065 5.270 1.735 ;
        RECT 3.145 0.610 3.595 0.940 ;
        RECT 3.765 0.895 4.775 1.065 ;
        RECT 3.765 0.440 3.935 0.895 ;
        RECT 2.805 0.270 3.935 0.440 ;
        RECT 4.105 0.085 4.435 0.725 ;
        RECT 4.605 0.425 4.775 0.895 ;
        RECT 4.945 0.595 5.275 1.065 ;
        RECT 5.445 1.010 5.615 1.820 ;
        RECT 6.285 1.630 6.455 2.240 ;
        RECT 6.625 1.970 6.955 2.980 ;
        RECT 7.125 2.140 7.455 3.245 ;
        RECT 8.235 2.140 8.485 3.245 ;
        RECT 6.625 1.800 7.535 1.970 ;
        RECT 9.155 1.820 9.485 3.245 ;
        RECT 7.365 1.630 7.535 1.800 ;
        RECT 6.285 1.300 7.030 1.630 ;
        RECT 7.365 1.300 8.435 1.630 ;
        RECT 7.365 1.130 7.535 1.300 ;
        RECT 5.445 0.425 5.835 1.010 ;
        RECT 4.605 0.255 5.835 0.425 ;
        RECT 6.005 0.085 6.335 1.010 ;
        RECT 6.825 0.960 7.535 1.130 ;
        RECT 6.825 0.350 7.155 0.960 ;
        RECT 7.385 0.085 7.635 0.790 ;
        RECT 8.295 0.085 8.545 0.790 ;
        RECT 9.235 0.085 9.485 1.130 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
  END
END sky130_fd_sc_hs__sdlclkp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__sedfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sedfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 6.575 1.180 7.075 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.060 0.835 1.780 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.450 2.085 1.780 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.075 1.180 5.635 1.510 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.450 4.865 1.780 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 16.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.190 1.175 8.160 1.240 ;
        RECT 4.300 1.140 8.160 1.175 ;
        RECT 14.655 1.140 16.315 1.260 ;
        RECT 4.300 1.115 12.730 1.140 ;
        RECT 1.600 1.000 12.730 1.115 ;
        RECT 0.005 0.920 12.730 1.000 ;
        RECT 13.700 0.920 16.315 1.140 ;
        RECT 0.005 0.245 16.315 0.920 ;
        RECT 0.000 0.000 16.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.510 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 16.320 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 14.845 1.820 15.240 2.980 ;
        RECT 14.845 0.620 15.015 1.820 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 15.860 1.820 16.235 2.980 ;
        RECT 16.065 1.150 16.235 1.820 ;
        RECT 15.875 0.370 16.235 1.150 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 16.320 3.415 ;
        RECT 0.115 2.460 0.445 2.980 ;
        RECT 0.955 2.630 1.205 3.245 ;
        RECT 1.375 2.905 2.225 3.075 ;
        RECT 1.375 2.460 1.545 2.905 ;
        RECT 0.115 2.290 1.545 2.460 ;
        RECT 0.115 0.810 0.285 2.290 ;
        RECT 1.715 2.120 1.885 2.735 ;
        RECT 2.055 2.480 2.225 2.905 ;
        RECT 2.395 2.650 2.645 3.245 ;
        RECT 3.185 2.480 3.545 2.980 ;
        RECT 2.055 2.310 3.545 2.480 ;
        RECT 1.025 1.950 2.665 2.120 ;
        RECT 1.025 1.280 1.355 1.950 ;
        RECT 2.335 1.525 2.665 1.950 ;
        RECT 2.875 1.525 3.205 2.140 ;
        RECT 3.375 1.345 3.545 2.310 ;
        RECT 1.025 1.110 2.040 1.280 ;
        RECT 0.115 0.480 0.660 0.810 ;
        RECT 1.150 0.085 1.480 0.890 ;
        RECT 1.710 0.545 2.040 1.110 ;
        RECT 3.030 1.175 3.545 1.345 ;
        RECT 3.715 2.905 4.785 3.075 ;
        RECT 3.715 2.300 3.965 2.905 ;
        RECT 2.210 0.085 2.540 1.005 ;
        RECT 3.030 0.545 3.360 1.175 ;
        RECT 3.715 1.005 3.885 2.300 ;
        RECT 4.135 2.290 4.445 2.735 ;
        RECT 4.615 2.460 4.785 2.905 ;
        RECT 4.955 2.630 5.205 3.245 ;
        RECT 5.715 2.480 6.045 2.970 ;
        RECT 6.275 2.650 6.605 3.245 ;
        RECT 7.665 2.650 7.995 3.245 ;
        RECT 8.165 2.730 9.020 2.980 ;
        RECT 8.165 2.480 8.335 2.730 ;
        RECT 9.190 2.560 9.520 2.980 ;
        RECT 10.080 2.730 10.410 3.245 ;
        RECT 11.175 2.730 11.505 3.245 ;
        RECT 5.715 2.460 8.335 2.480 ;
        RECT 4.615 2.310 8.335 2.460 ;
        RECT 9.040 2.390 9.520 2.560 ;
        RECT 9.690 2.390 12.595 2.560 ;
        RECT 12.765 2.520 13.195 2.980 ;
        RECT 13.640 2.650 14.230 3.245 ;
        RECT 4.615 2.290 6.210 2.310 ;
        RECT 4.135 2.120 4.305 2.290 ;
        RECT 3.530 0.545 3.885 1.005 ;
        RECT 4.055 1.950 5.870 2.120 ;
        RECT 4.055 1.065 4.305 1.950 ;
        RECT 5.565 1.790 5.870 1.950 ;
        RECT 4.055 0.605 4.740 1.065 ;
        RECT 6.040 1.010 6.210 2.290 ;
        RECT 6.725 1.820 7.525 2.140 ;
        RECT 7.055 1.810 7.525 1.820 ;
        RECT 7.355 1.010 7.525 1.810 ;
        RECT 7.775 1.650 7.945 2.310 ;
        RECT 8.585 2.140 8.870 2.380 ;
        RECT 8.115 1.820 8.870 2.140 ;
        RECT 7.775 1.480 8.530 1.650 ;
        RECT 4.055 0.410 4.305 0.605 ;
        RECT 4.910 0.085 5.240 1.010 ;
        RECT 5.740 0.605 6.210 1.010 ;
        RECT 6.380 0.085 6.550 1.010 ;
        RECT 6.730 0.840 7.525 1.010 ;
        RECT 6.730 0.350 7.060 0.840 ;
        RECT 7.290 0.085 7.620 0.670 ;
        RECT 7.800 0.425 8.050 1.130 ;
        RECT 8.280 0.595 8.530 1.480 ;
        RECT 8.700 0.425 8.870 1.820 ;
        RECT 9.040 1.790 9.210 2.390 ;
        RECT 9.690 2.220 9.860 2.390 ;
        RECT 9.380 1.960 9.860 2.220 ;
        RECT 10.615 2.050 11.070 2.220 ;
        RECT 10.400 1.790 10.730 1.830 ;
        RECT 9.040 1.620 10.730 1.790 ;
        RECT 9.040 0.950 9.210 1.620 ;
        RECT 10.400 1.530 10.730 1.620 ;
        RECT 10.900 1.520 11.070 2.050 ;
        RECT 12.425 1.800 12.595 2.390 ;
        RECT 13.025 1.885 13.195 2.520 ;
        RECT 14.430 2.380 14.600 2.980 ;
        RECT 13.460 2.055 14.600 2.380 ;
        RECT 14.045 1.920 14.600 2.055 ;
        RECT 9.380 1.120 9.690 1.450 ;
        RECT 9.860 1.360 10.190 1.450 ;
        RECT 10.900 1.360 11.740 1.520 ;
        RECT 9.860 1.190 11.740 1.360 ;
        RECT 11.950 1.300 12.255 1.800 ;
        RECT 12.425 1.470 12.855 1.800 ;
        RECT 13.025 1.715 13.875 1.885 ;
        RECT 13.065 1.300 13.395 1.545 ;
        RECT 9.490 1.020 9.690 1.120 ;
        RECT 9.040 0.620 9.320 0.950 ;
        RECT 9.490 0.850 10.730 1.020 ;
        RECT 9.490 0.425 9.690 0.850 ;
        RECT 7.800 0.255 9.690 0.425 ;
        RECT 10.065 0.085 10.390 0.680 ;
        RECT 10.560 0.425 10.730 0.850 ;
        RECT 10.900 0.595 11.070 1.190 ;
        RECT 11.950 1.130 13.395 1.300 ;
        RECT 13.705 1.530 13.875 1.715 ;
        RECT 13.705 1.200 14.260 1.530 ;
        RECT 11.950 1.020 12.120 1.130 ;
        RECT 11.240 0.850 12.120 1.020 ;
        RECT 13.705 0.940 13.875 1.200 ;
        RECT 14.430 1.030 14.600 1.920 ;
        RECT 15.440 1.820 15.690 3.245 ;
        RECT 11.240 0.425 11.410 0.850 ;
        RECT 12.290 0.770 13.875 0.940 ;
        RECT 10.560 0.255 11.410 0.425 ;
        RECT 11.580 0.085 11.830 0.680 ;
        RECT 12.290 0.350 12.620 0.770 ;
        RECT 13.190 0.085 14.035 0.600 ;
        RECT 14.205 0.425 14.600 1.030 ;
        RECT 15.185 1.320 15.895 1.650 ;
        RECT 15.185 0.425 15.355 1.320 ;
        RECT 14.205 0.255 15.355 0.425 ;
        RECT 15.525 0.085 15.695 1.150 ;
        RECT 0.000 -0.085 16.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 3.035 1.950 3.205 2.120 ;
        RECT 14.075 1.950 14.245 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
      LAYER met1 ;
        RECT 2.975 2.105 3.265 2.150 ;
        RECT 14.015 2.105 14.305 2.150 ;
        RECT 2.975 1.965 14.305 2.105 ;
        RECT 2.975 1.920 3.265 1.965 ;
        RECT 14.015 1.920 14.305 1.965 ;
  END
END sky130_fd_sc_hs__sedfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sedfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 6.705 1.180 7.045 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.980 0.835 1.990 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.450 1.905 1.780 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.125 1.180 5.635 1.510 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.180 4.915 1.510 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 17.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.305 1.175 8.345 1.240 ;
        RECT 4.350 1.115 8.345 1.175 ;
        RECT 1.570 1.035 8.345 1.115 ;
        RECT 10.445 1.035 12.860 1.140 ;
        RECT 1.570 0.920 12.860 1.035 ;
        RECT 13.885 0.920 17.225 1.240 ;
        RECT 0.030 0.245 17.225 0.920 ;
        RECT 0.000 0.000 17.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 17.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 17.280 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 15.485 0.350 15.825 2.150 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 16.435 1.975 16.665 3.010 ;
        RECT 16.435 1.805 17.165 1.975 ;
        RECT 16.700 1.130 17.165 1.805 ;
        RECT 16.355 0.960 17.165 1.130 ;
        RECT 16.355 0.350 16.685 0.960 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 17.280 3.415 ;
        RECT 0.085 2.460 0.525 2.980 ;
        RECT 1.065 2.630 1.315 3.245 ;
        RECT 1.485 2.905 2.335 3.075 ;
        RECT 1.485 2.460 1.655 2.905 ;
        RECT 0.085 2.290 1.655 2.460 ;
        RECT 0.085 0.730 0.255 2.290 ;
        RECT 1.825 2.120 1.995 2.735 ;
        RECT 2.165 2.460 2.335 2.905 ;
        RECT 2.505 2.630 2.755 3.245 ;
        RECT 3.265 2.460 3.545 2.970 ;
        RECT 2.165 2.290 3.545 2.460 ;
        RECT 1.005 1.950 2.635 2.120 ;
        RECT 1.005 1.280 1.335 1.950 ;
        RECT 2.305 1.515 2.635 1.950 ;
        RECT 2.875 1.515 3.205 1.845 ;
        RECT 3.375 1.345 3.545 2.290 ;
        RECT 1.005 1.110 2.010 1.280 ;
        RECT 0.085 0.420 0.580 0.730 ;
        RECT 1.070 0.085 1.400 0.810 ;
        RECT 1.680 0.545 2.010 1.110 ;
        RECT 3.000 1.175 3.545 1.345 ;
        RECT 3.715 2.905 4.865 3.075 ;
        RECT 3.715 2.290 3.965 2.905 ;
        RECT 2.180 0.085 2.510 1.005 ;
        RECT 3.000 0.545 3.330 1.175 ;
        RECT 3.715 1.005 3.885 2.290 ;
        RECT 4.135 2.245 4.525 2.735 ;
        RECT 4.695 2.425 4.865 2.905 ;
        RECT 5.035 2.595 5.305 3.245 ;
        RECT 5.845 2.480 6.305 2.925 ;
        RECT 6.485 2.650 6.735 3.245 ;
        RECT 7.795 2.650 8.125 3.245 ;
        RECT 8.805 2.650 9.055 2.980 ;
        RECT 8.295 2.480 9.055 2.650 ;
        RECT 9.225 2.530 9.585 2.980 ;
        RECT 10.225 2.730 10.555 3.245 ;
        RECT 11.320 2.730 11.650 3.245 ;
        RECT 5.845 2.425 8.465 2.480 ;
        RECT 4.695 2.310 8.465 2.425 ;
        RECT 4.695 2.255 6.475 2.310 ;
        RECT 4.135 2.055 4.305 2.245 ;
        RECT 3.500 0.545 3.885 1.005 ;
        RECT 4.055 1.850 4.305 2.055 ;
        RECT 5.805 1.850 6.135 2.085 ;
        RECT 4.055 1.680 6.135 1.850 ;
        RECT 4.055 1.010 4.305 1.680 ;
        RECT 5.805 1.430 6.135 1.680 ;
        RECT 6.305 1.260 6.475 2.255 ;
        RECT 6.855 1.820 7.655 2.140 ;
        RECT 5.820 1.090 6.475 1.260 ;
        RECT 7.215 1.470 7.655 1.820 ;
        RECT 7.905 1.650 8.075 2.310 ;
        RECT 8.725 2.140 9.055 2.305 ;
        RECT 8.245 1.820 9.055 2.140 ;
        RECT 7.905 1.480 8.715 1.650 ;
        RECT 4.055 0.605 4.790 1.010 ;
        RECT 4.055 0.365 4.305 0.605 ;
        RECT 4.960 0.085 5.290 1.010 ;
        RECT 5.820 0.605 6.150 1.090 ;
        RECT 7.215 1.010 7.385 1.470 ;
        RECT 6.415 0.085 6.745 0.920 ;
        RECT 6.915 0.350 7.385 1.010 ;
        RECT 7.555 0.085 7.725 1.130 ;
        RECT 7.905 0.425 8.235 1.130 ;
        RECT 8.465 0.595 8.715 1.480 ;
        RECT 8.885 0.425 9.055 1.820 ;
        RECT 9.225 1.860 9.395 2.530 ;
        RECT 9.755 2.390 12.720 2.560 ;
        RECT 12.890 2.520 13.325 2.980 ;
        RECT 13.765 2.650 14.305 3.245 ;
        RECT 9.755 2.360 9.925 2.390 ;
        RECT 9.565 2.030 9.925 2.360 ;
        RECT 10.760 2.050 11.385 2.220 ;
        RECT 9.225 1.690 10.940 1.860 ;
        RECT 9.225 0.595 9.395 1.690 ;
        RECT 10.610 1.530 10.940 1.690 ;
        RECT 11.215 1.520 11.385 2.050 ;
        RECT 12.550 1.800 12.720 2.390 ;
        RECT 13.155 1.885 13.325 2.520 ;
        RECT 14.475 2.490 14.835 2.980 ;
        RECT 15.035 2.660 15.365 3.245 ;
        RECT 15.935 2.660 16.265 3.245 ;
        RECT 14.475 2.380 16.185 2.490 ;
        RECT 13.585 2.320 16.185 2.380 ;
        RECT 13.585 2.055 15.235 2.320 ;
        RECT 10.065 1.360 10.395 1.520 ;
        RECT 11.215 1.360 11.885 1.520 ;
        RECT 9.565 1.020 9.855 1.345 ;
        RECT 10.065 1.190 11.885 1.360 ;
        RECT 12.080 1.300 12.380 1.800 ;
        RECT 12.550 1.470 12.985 1.800 ;
        RECT 13.155 1.715 13.865 1.885 ;
        RECT 14.475 1.800 15.235 2.055 ;
        RECT 13.695 1.630 13.865 1.715 ;
        RECT 13.195 1.300 13.525 1.545 ;
        RECT 9.565 0.850 10.860 1.020 ;
        RECT 9.565 0.425 9.735 0.850 ;
        RECT 7.905 0.255 9.735 0.425 ;
        RECT 10.270 0.085 10.520 0.680 ;
        RECT 10.690 0.425 10.860 0.850 ;
        RECT 11.030 0.595 11.200 1.190 ;
        RECT 12.080 1.130 13.525 1.300 ;
        RECT 13.695 1.300 14.495 1.630 ;
        RECT 14.665 1.550 15.235 1.800 ;
        RECT 15.995 1.635 16.185 2.320 ;
        RECT 16.835 2.145 17.165 3.245 ;
        RECT 12.080 1.020 12.250 1.130 ;
        RECT 11.370 0.850 12.250 1.020 ;
        RECT 13.695 0.940 13.865 1.300 ;
        RECT 14.665 1.130 14.835 1.550 ;
        RECT 15.995 1.300 16.510 1.635 ;
        RECT 11.370 0.425 11.540 0.850 ;
        RECT 12.420 0.770 13.865 0.940 ;
        RECT 10.690 0.255 11.540 0.425 ;
        RECT 11.710 0.085 11.960 0.680 ;
        RECT 12.420 0.350 12.750 0.770 ;
        RECT 14.065 0.600 14.335 1.120 ;
        RECT 13.320 0.085 14.335 0.600 ;
        RECT 14.505 0.350 14.835 1.130 ;
        RECT 15.065 0.085 15.315 1.130 ;
        RECT 16.005 0.085 16.175 1.130 ;
        RECT 16.855 0.085 17.115 0.790 ;
        RECT 0.000 -0.085 17.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 16.955 3.245 17.125 3.415 ;
        RECT 3.035 1.580 3.205 1.750 ;
        RECT 15.035 1.580 15.205 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
        RECT 16.955 -0.085 17.125 0.085 ;
      LAYER met1 ;
        RECT 2.975 1.735 3.265 1.780 ;
        RECT 14.975 1.735 15.265 1.780 ;
        RECT 2.975 1.595 15.265 1.735 ;
        RECT 2.975 1.550 3.265 1.595 ;
        RECT 14.975 1.550 15.265 1.595 ;
  END
END sky130_fd_sc_hs__sedfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sedfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sedfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 6.330 1.180 6.660 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.110 0.805 1.780 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.320 1.845 1.780 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.180 5.280 1.745 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.400 1.180 4.730 1.510 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 15.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.910 1.175 7.870 1.240 ;
        RECT 4.140 1.105 7.870 1.175 ;
        RECT 1.530 1.035 7.870 1.105 ;
        RECT 9.925 1.035 12.340 1.140 ;
        RECT 1.530 0.920 12.340 1.035 ;
        RECT 14.375 0.920 15.355 1.240 ;
        RECT 0.005 0.245 15.355 0.920 ;
        RECT 0.000 0.000 15.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 15.550 3.520 ;
        RECT 6.020 1.600 7.080 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 15.360 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.518900 ;
    PORT
      LAYER li1 ;
        RECT 14.475 0.350 14.815 2.980 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 15.360 3.415 ;
        RECT 0.085 2.460 0.435 2.980 ;
        RECT 0.945 2.630 1.195 3.245 ;
        RECT 1.365 2.905 2.215 3.075 ;
        RECT 1.365 2.460 1.535 2.905 ;
        RECT 0.085 2.290 1.535 2.460 ;
        RECT 0.085 0.810 0.255 2.290 ;
        RECT 1.705 2.120 1.875 2.735 ;
        RECT 2.045 2.460 2.215 2.905 ;
        RECT 2.385 2.630 2.635 3.245 ;
        RECT 3.145 2.460 3.395 2.975 ;
        RECT 2.045 2.290 3.395 2.460 ;
        RECT 0.975 1.950 2.385 2.120 ;
        RECT 0.975 1.150 1.305 1.950 ;
        RECT 2.055 1.520 2.385 1.950 ;
        RECT 2.555 1.505 3.055 1.835 ;
        RECT 3.225 1.335 3.395 2.290 ;
        RECT 2.890 1.165 3.395 1.335 ;
        RECT 3.565 2.905 4.710 3.075 ;
        RECT 3.565 2.295 3.845 2.905 ;
        RECT 0.975 0.995 1.810 1.150 ;
        RECT 0.975 0.980 1.890 0.995 ;
        RECT 0.085 0.480 0.590 0.810 ;
        RECT 1.080 0.085 1.410 0.810 ;
        RECT 1.640 0.535 1.890 0.980 ;
        RECT 2.070 0.085 2.400 0.995 ;
        RECT 2.890 0.535 3.220 1.165 ;
        RECT 3.565 0.995 3.735 2.295 ;
        RECT 4.015 2.255 4.370 2.735 ;
        RECT 4.540 2.425 4.710 2.905 ;
        RECT 4.880 2.595 5.130 3.245 ;
        RECT 5.640 2.500 5.990 2.935 ;
        RECT 6.160 2.670 6.490 3.245 ;
        RECT 7.510 2.670 7.840 3.245 ;
        RECT 8.010 2.730 8.815 2.980 ;
        RECT 8.010 2.500 8.180 2.730 ;
        RECT 8.985 2.560 9.315 2.980 ;
        RECT 9.865 2.730 10.195 3.245 ;
        RECT 10.905 2.730 11.235 3.245 ;
        RECT 5.640 2.425 8.180 2.500 ;
        RECT 4.540 2.330 8.180 2.425 ;
        RECT 8.835 2.390 9.315 2.560 ;
        RECT 9.485 2.390 12.200 2.560 ;
        RECT 4.540 2.255 6.160 2.330 ;
        RECT 4.015 2.085 4.185 2.255 ;
        RECT 3.390 0.535 3.735 0.995 ;
        RECT 3.905 1.915 5.820 2.085 ;
        RECT 3.905 1.010 4.185 1.915 ;
        RECT 5.490 1.415 5.820 1.915 ;
        RECT 5.990 1.245 6.160 2.255 ;
        RECT 6.610 1.830 7.390 2.160 ;
        RECT 6.610 1.760 7.000 1.830 ;
        RECT 5.465 1.075 6.160 1.245 ;
        RECT 3.905 0.605 4.575 1.010 ;
        RECT 3.905 0.255 4.185 0.605 ;
        RECT 4.755 0.085 5.005 1.010 ;
        RECT 5.465 0.605 5.795 1.075 ;
        RECT 6.830 1.010 7.000 1.760 ;
        RECT 7.620 1.650 7.790 2.330 ;
        RECT 8.405 2.160 8.665 2.335 ;
        RECT 7.960 1.990 8.665 2.160 ;
        RECT 7.960 1.820 8.575 1.990 ;
        RECT 7.620 1.480 8.235 1.650 ;
        RECT 6.020 0.085 6.280 0.905 ;
        RECT 6.450 0.840 7.000 1.010 ;
        RECT 6.450 0.350 6.780 0.840 ;
        RECT 7.005 0.085 7.335 0.670 ;
        RECT 7.515 0.425 7.765 1.130 ;
        RECT 7.985 0.595 8.235 1.480 ;
        RECT 8.405 0.425 8.575 1.820 ;
        RECT 8.835 1.790 9.005 2.390 ;
        RECT 9.485 2.220 9.655 2.390 ;
        RECT 9.175 1.960 9.655 2.220 ;
        RECT 10.385 1.970 10.805 2.220 ;
        RECT 10.135 1.790 10.465 1.795 ;
        RECT 8.745 1.620 10.465 1.790 ;
        RECT 8.745 0.595 8.915 1.620 ;
        RECT 10.135 1.535 10.465 1.620 ;
        RECT 10.635 1.525 10.805 1.970 ;
        RECT 9.565 1.365 9.895 1.450 ;
        RECT 10.635 1.365 11.385 1.525 ;
        RECT 9.085 1.020 9.340 1.345 ;
        RECT 9.565 1.195 11.385 1.365 ;
        RECT 11.560 1.280 11.860 1.800 ;
        RECT 12.030 1.735 12.200 2.390 ;
        RECT 12.370 1.940 12.805 2.980 ;
        RECT 13.330 2.650 13.785 3.245 ;
        RECT 13.955 2.380 14.285 2.980 ;
        RECT 13.065 2.075 14.285 2.380 ;
        RECT 12.635 1.905 12.805 1.940 ;
        RECT 12.635 1.735 13.785 1.905 ;
        RECT 12.030 1.450 12.465 1.735 ;
        RECT 12.675 1.280 13.005 1.555 ;
        RECT 9.565 1.190 9.895 1.195 ;
        RECT 9.085 0.850 10.340 1.020 ;
        RECT 9.085 0.425 9.255 0.850 ;
        RECT 7.515 0.255 9.255 0.425 ;
        RECT 9.750 0.085 10.000 0.680 ;
        RECT 10.170 0.425 10.340 0.850 ;
        RECT 10.510 0.595 10.680 1.195 ;
        RECT 11.560 1.110 13.005 1.280 ;
        RECT 11.560 1.025 11.730 1.110 ;
        RECT 10.850 0.855 11.730 1.025 ;
        RECT 13.175 0.940 13.345 1.735 ;
        RECT 13.615 1.380 13.785 1.735 ;
        RECT 14.045 1.550 14.285 2.075 ;
        RECT 15.005 1.820 15.255 3.245 ;
        RECT 13.615 1.050 13.945 1.380 ;
        RECT 10.850 0.425 11.020 0.855 ;
        RECT 11.900 0.770 13.345 0.940 ;
        RECT 14.115 0.810 14.285 1.550 ;
        RECT 10.170 0.255 11.020 0.425 ;
        RECT 11.190 0.085 11.440 0.685 ;
        RECT 11.900 0.350 12.230 0.770 ;
        RECT 12.800 0.085 13.755 0.600 ;
        RECT 13.925 0.350 14.285 0.810 ;
        RECT 14.995 0.085 15.245 1.130 ;
        RECT 0.000 -0.085 15.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 2.555 1.580 2.725 1.750 ;
        RECT 14.075 1.580 14.245 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
      LAYER met1 ;
        RECT 2.495 1.735 2.785 1.780 ;
        RECT 14.015 1.735 14.305 1.780 ;
        RECT 2.495 1.595 14.305 1.735 ;
        RECT 2.495 1.550 2.785 1.595 ;
        RECT 14.015 1.550 14.305 1.595 ;
  END
END sky130_fd_sc_hs__sedfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hs__sedfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sedfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 6.395 1.180 6.725 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.980 0.805 1.990 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.320 1.845 1.780 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 4.955 1.180 5.410 1.745 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.465 1.180 4.785 1.510 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 16.320 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.125 1.175 8.105 1.240 ;
        RECT 4.275 1.115 8.105 1.175 ;
        RECT 1.505 1.035 8.105 1.115 ;
        RECT 10.290 1.035 12.750 1.140 ;
        RECT 1.505 0.920 12.750 1.035 ;
        RECT 14.765 0.920 16.315 1.240 ;
        RECT 0.125 0.245 16.315 0.920 ;
        RECT 0.000 0.000 16.320 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.510 3.520 ;
        RECT 6.200 1.640 7.305 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 16.320 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.560000 ;
    PORT
      LAYER li1 ;
        RECT 15.460 2.150 15.705 2.980 ;
        RECT 15.460 1.550 16.195 2.150 ;
        RECT 15.460 1.130 15.705 1.550 ;
        RECT 15.375 0.350 15.705 1.130 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 16.320 3.415 ;
        RECT 0.085 2.460 0.510 2.980 ;
        RECT 1.050 2.630 1.300 3.245 ;
        RECT 1.470 2.905 2.320 3.075 ;
        RECT 1.470 2.460 1.640 2.905 ;
        RECT 0.085 2.290 1.640 2.460 ;
        RECT 0.085 0.810 0.255 2.290 ;
        RECT 1.810 2.120 1.980 2.735 ;
        RECT 2.150 2.460 2.320 2.905 ;
        RECT 2.490 2.630 2.740 3.245 ;
        RECT 3.250 2.460 3.500 2.975 ;
        RECT 2.150 2.290 3.500 2.460 ;
        RECT 0.975 1.950 2.385 2.120 ;
        RECT 0.975 1.150 1.305 1.950 ;
        RECT 2.055 1.520 2.385 1.950 ;
        RECT 2.555 1.515 3.070 1.845 ;
        RECT 3.330 1.345 3.500 2.290 ;
        RECT 3.170 1.175 3.500 1.345 ;
        RECT 3.670 2.905 4.840 3.075 ;
        RECT 3.670 2.295 3.950 2.905 ;
        RECT 0.975 0.980 1.865 1.150 ;
        RECT 3.170 1.005 3.340 1.175 ;
        RECT 3.670 1.005 3.840 2.295 ;
        RECT 4.125 2.255 4.500 2.735 ;
        RECT 4.670 2.425 4.840 2.905 ;
        RECT 5.010 2.595 5.260 3.245 ;
        RECT 5.800 2.540 6.130 2.935 ;
        RECT 6.360 2.710 6.695 3.245 ;
        RECT 7.755 2.710 8.085 3.245 ;
        RECT 8.765 2.690 9.015 2.980 ;
        RECT 8.255 2.540 9.015 2.690 ;
        RECT 5.800 2.520 9.015 2.540 ;
        RECT 9.185 2.520 9.545 2.980 ;
        RECT 10.215 2.730 10.545 3.245 ;
        RECT 11.310 2.730 11.650 3.245 ;
        RECT 5.800 2.425 8.425 2.520 ;
        RECT 4.670 2.370 8.425 2.425 ;
        RECT 4.670 2.255 6.225 2.370 ;
        RECT 4.125 2.085 4.295 2.255 ;
        RECT 0.085 0.350 0.565 0.810 ;
        RECT 1.055 0.085 1.385 0.810 ;
        RECT 1.615 0.545 1.865 0.980 ;
        RECT 2.045 0.085 2.375 1.005 ;
        RECT 2.865 0.675 3.340 1.005 ;
        RECT 3.510 0.545 3.840 1.005 ;
        RECT 4.010 1.915 5.885 2.085 ;
        RECT 4.010 1.010 4.295 1.915 ;
        RECT 5.620 1.415 5.885 1.915 ;
        RECT 6.055 1.065 6.225 2.255 ;
        RECT 4.010 0.605 4.715 1.010 ;
        RECT 4.010 0.255 4.295 0.605 ;
        RECT 4.885 0.085 5.215 1.010 ;
        RECT 5.675 0.895 6.225 1.065 ;
        RECT 6.895 1.530 7.615 2.200 ;
        RECT 7.865 1.650 8.035 2.370 ;
        RECT 8.645 2.200 9.005 2.350 ;
        RECT 8.205 2.020 9.005 2.200 ;
        RECT 8.205 1.820 8.815 2.020 ;
        RECT 9.185 1.830 9.355 2.520 ;
        RECT 9.715 2.390 12.730 2.560 ;
        RECT 9.715 2.350 9.885 2.390 ;
        RECT 9.525 2.020 9.885 2.350 ;
        RECT 10.750 2.050 11.125 2.220 ;
        RECT 6.895 1.010 7.065 1.530 ;
        RECT 7.865 1.480 8.475 1.650 ;
        RECT 5.675 0.605 6.005 0.895 ;
        RECT 6.235 0.085 6.495 0.680 ;
        RECT 6.675 0.350 7.065 1.010 ;
        RECT 7.235 0.085 7.485 1.130 ;
        RECT 7.665 0.425 7.995 1.130 ;
        RECT 8.225 0.595 8.475 1.480 ;
        RECT 8.645 0.425 8.815 1.820 ;
        RECT 8.985 1.660 10.785 1.830 ;
        RECT 8.985 0.595 9.155 1.660 ;
        RECT 10.455 1.530 10.785 1.660 ;
        RECT 10.955 1.520 11.125 2.050 ;
        RECT 9.915 1.360 10.245 1.490 ;
        RECT 10.955 1.360 11.800 1.520 ;
        RECT 9.325 1.020 9.655 1.345 ;
        RECT 9.915 1.190 11.800 1.360 ;
        RECT 12.040 1.360 12.370 1.800 ;
        RECT 12.560 1.755 12.730 2.390 ;
        RECT 12.900 1.925 13.250 2.980 ;
        RECT 13.690 2.650 14.230 3.245 ;
        RECT 14.400 2.470 14.750 2.980 ;
        RECT 13.510 2.300 14.750 2.470 ;
        RECT 13.510 2.095 13.840 2.300 ;
        RECT 14.080 1.925 14.410 2.130 ;
        RECT 13.080 1.755 14.410 1.925 ;
        RECT 12.560 1.530 12.910 1.755 ;
        RECT 13.120 1.360 13.450 1.585 ;
        RECT 12.040 1.190 13.450 1.360 ;
        RECT 9.325 0.850 10.705 1.020 ;
        RECT 9.325 0.425 9.495 0.850 ;
        RECT 7.665 0.255 9.495 0.425 ;
        RECT 10.100 0.085 10.365 0.680 ;
        RECT 10.535 0.425 10.705 0.850 ;
        RECT 10.875 0.595 11.125 1.190 ;
        RECT 12.040 1.020 12.210 1.190 ;
        RECT 13.620 1.020 13.790 1.755 ;
        RECT 14.080 1.460 14.410 1.755 ;
        RECT 14.580 1.780 14.750 2.300 ;
        RECT 14.960 1.950 15.290 3.245 ;
        RECT 15.875 2.320 16.205 3.245 ;
        RECT 14.580 1.550 15.235 1.780 ;
        RECT 14.580 1.290 14.750 1.550 ;
        RECT 11.295 0.850 12.210 1.020 ;
        RECT 12.390 0.850 13.790 1.020 ;
        RECT 14.315 1.120 14.750 1.290 ;
        RECT 11.295 0.425 11.465 0.850 ;
        RECT 10.535 0.255 11.465 0.425 ;
        RECT 11.635 0.085 11.885 0.680 ;
        RECT 12.390 0.350 12.720 0.850 ;
        RECT 13.210 0.085 14.145 0.680 ;
        RECT 14.315 0.350 14.645 1.120 ;
        RECT 14.875 0.085 15.205 0.950 ;
        RECT 15.875 0.085 16.205 1.130 ;
        RECT 0.000 -0.085 16.320 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 2.555 1.580 2.725 1.750 ;
        RECT 15.035 1.580 15.205 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
      LAYER met1 ;
        RECT 2.495 1.735 2.785 1.780 ;
        RECT 14.975 1.735 15.265 1.780 ;
        RECT 2.495 1.595 15.265 1.735 ;
        RECT 2.495 1.550 2.785 1.595 ;
        RECT 14.975 1.550 15.265 1.595 ;
  END
END sky130_fd_sc_hs__sedfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hs__sedfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sedfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 6.455 1.180 7.075 1.550 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.980 0.825 1.990 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.320 1.865 1.780 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 4.955 1.180 5.370 1.745 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.180 4.785 1.510 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 16.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.000 1.175 7.960 1.240 ;
        RECT 4.225 1.115 7.960 1.175 ;
        RECT 1.490 1.035 7.960 1.115 ;
        RECT 10.015 1.140 10.960 1.165 ;
        RECT 10.015 1.035 12.395 1.140 ;
        RECT 1.490 0.920 12.395 1.035 ;
        RECT 14.455 0.920 16.795 1.450 ;
        RECT 0.110 0.245 16.795 0.920 ;
        RECT 0.000 0.000 16.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 16.990 3.520 ;
        RECT 6.115 1.625 7.180 1.660 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 16.800 3.575 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.097500 ;
    PORT
      LAYER li1 ;
        RECT 15.065 2.150 15.285 2.980 ;
        RECT 15.970 2.150 16.185 2.980 ;
        RECT 15.065 1.820 16.675 2.150 ;
        RECT 15.165 1.340 16.675 1.820 ;
        RECT 15.075 1.090 16.675 1.340 ;
        RECT 15.075 0.560 15.325 1.090 ;
        RECT 15.995 0.575 16.200 1.090 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 16.800 3.415 ;
        RECT 0.085 2.460 0.495 2.980 ;
        RECT 1.035 2.630 1.285 3.245 ;
        RECT 1.455 2.905 2.305 3.075 ;
        RECT 1.455 2.460 1.625 2.905 ;
        RECT 0.085 2.290 1.625 2.460 ;
        RECT 0.085 0.810 0.255 2.290 ;
        RECT 1.795 2.120 1.965 2.735 ;
        RECT 2.135 2.460 2.305 2.905 ;
        RECT 2.475 2.630 2.725 3.245 ;
        RECT 3.235 2.460 3.485 2.975 ;
        RECT 2.135 2.290 3.485 2.460 ;
        RECT 0.995 1.950 2.365 2.120 ;
        RECT 0.995 1.150 1.325 1.950 ;
        RECT 2.115 1.520 2.365 1.950 ;
        RECT 2.535 1.520 3.055 1.850 ;
        RECT 3.315 1.345 3.485 2.290 ;
        RECT 2.850 1.175 3.485 1.345 ;
        RECT 3.655 2.905 4.800 3.075 ;
        RECT 3.655 2.295 3.935 2.905 ;
        RECT 0.995 0.980 1.850 1.150 ;
        RECT 0.085 0.340 0.550 0.810 ;
        RECT 1.040 0.085 1.370 0.810 ;
        RECT 1.600 0.545 1.850 0.980 ;
        RECT 2.030 0.085 2.360 1.005 ;
        RECT 2.850 0.545 3.180 1.175 ;
        RECT 3.655 1.005 3.825 2.295 ;
        RECT 4.105 2.255 4.460 2.735 ;
        RECT 4.630 2.425 4.800 2.905 ;
        RECT 4.970 2.595 5.220 3.245 ;
        RECT 5.730 2.505 6.060 2.935 ;
        RECT 6.260 2.675 6.590 3.245 ;
        RECT 7.610 2.675 7.940 3.245 ;
        RECT 8.155 2.505 8.830 2.980 ;
        RECT 9.000 2.520 9.360 2.980 ;
        RECT 9.960 2.730 10.290 3.245 ;
        RECT 10.995 2.730 11.325 3.245 ;
        RECT 5.730 2.425 8.325 2.505 ;
        RECT 4.630 2.335 8.325 2.425 ;
        RECT 4.630 2.255 6.200 2.335 ;
        RECT 4.105 2.085 4.275 2.255 ;
        RECT 3.350 0.675 3.825 1.005 ;
        RECT 3.995 1.915 5.860 2.085 ;
        RECT 3.995 1.010 4.275 1.915 ;
        RECT 5.580 1.415 5.860 1.915 ;
        RECT 6.030 1.245 6.200 2.255 ;
        RECT 6.710 1.785 7.490 2.165 ;
        RECT 5.555 1.075 6.200 1.245 ;
        RECT 3.995 0.605 4.585 1.010 ;
        RECT 3.995 0.255 4.275 0.605 ;
        RECT 4.765 0.085 5.095 1.010 ;
        RECT 5.555 0.605 5.885 1.075 ;
        RECT 7.245 1.010 7.415 1.785 ;
        RECT 7.720 1.650 7.890 2.335 ;
        RECT 8.495 2.165 8.830 2.335 ;
        RECT 8.060 1.995 8.830 2.165 ;
        RECT 8.060 1.820 8.665 1.995 ;
        RECT 7.720 1.480 8.325 1.650 ;
        RECT 6.110 0.085 6.360 0.905 ;
        RECT 6.540 0.840 7.415 1.010 ;
        RECT 6.540 0.350 6.870 0.840 ;
        RECT 7.095 0.085 7.425 0.670 ;
        RECT 7.605 0.425 7.855 1.130 ;
        RECT 8.075 0.595 8.325 1.480 ;
        RECT 8.495 0.425 8.665 1.820 ;
        RECT 9.000 1.800 9.170 2.520 ;
        RECT 9.530 2.390 12.295 2.560 ;
        RECT 9.530 2.330 9.700 2.390 ;
        RECT 9.340 2.000 9.700 2.330 ;
        RECT 10.475 1.970 10.925 2.220 ;
        RECT 8.835 1.630 10.585 1.800 ;
        RECT 8.835 0.595 9.005 1.630 ;
        RECT 10.255 1.540 10.585 1.630 ;
        RECT 10.755 1.530 10.925 1.970 ;
        RECT 9.715 1.370 10.045 1.405 ;
        RECT 10.755 1.370 11.475 1.530 ;
        RECT 9.175 1.030 9.505 1.255 ;
        RECT 9.715 1.200 11.475 1.370 ;
        RECT 11.685 1.360 11.955 1.800 ;
        RECT 12.125 1.755 12.295 2.390 ;
        RECT 12.465 1.925 12.895 2.980 ;
        RECT 13.335 2.650 13.875 3.245 ;
        RECT 14.045 2.350 14.395 2.980 ;
        RECT 13.155 2.180 14.395 2.350 ;
        RECT 13.155 2.095 13.485 2.180 ;
        RECT 13.725 1.925 14.055 1.990 ;
        RECT 12.725 1.755 14.055 1.925 ;
        RECT 12.125 1.530 12.555 1.755 ;
        RECT 12.765 1.360 13.095 1.585 ;
        RECT 9.175 0.860 10.430 1.030 ;
        RECT 9.175 0.425 9.505 0.860 ;
        RECT 7.605 0.255 9.505 0.425 ;
        RECT 9.840 0.085 10.090 0.690 ;
        RECT 10.260 0.425 10.430 0.860 ;
        RECT 10.600 0.595 10.770 1.200 ;
        RECT 11.685 1.190 13.095 1.360 ;
        RECT 11.685 1.030 11.855 1.190 ;
        RECT 10.940 0.860 11.855 1.030 ;
        RECT 13.265 1.020 14.055 1.755 ;
        RECT 12.035 0.990 14.055 1.020 ;
        RECT 10.940 0.425 11.110 0.860 ;
        RECT 12.035 0.850 13.435 0.990 ;
        RECT 13.725 0.980 14.055 0.990 ;
        RECT 14.225 1.780 14.395 2.180 ;
        RECT 14.565 1.950 14.895 3.245 ;
        RECT 15.465 2.320 15.795 3.245 ;
        RECT 16.365 2.320 16.695 3.245 ;
        RECT 14.225 1.550 14.755 1.780 ;
        RECT 10.260 0.255 11.110 0.425 ;
        RECT 11.280 0.085 11.530 0.690 ;
        RECT 12.035 0.350 12.365 0.850 ;
        RECT 14.225 0.810 14.395 1.550 ;
        RECT 12.855 0.085 13.835 0.680 ;
        RECT 14.005 0.350 14.395 0.810 ;
        RECT 14.565 0.085 14.895 1.340 ;
        RECT 15.495 0.085 15.825 0.920 ;
        RECT 16.370 0.085 16.700 0.920 ;
        RECT 0.000 -0.085 16.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 15.515 3.245 15.685 3.415 ;
        RECT 15.995 3.245 16.165 3.415 ;
        RECT 16.475 3.245 16.645 3.415 ;
        RECT 2.555 1.580 2.725 1.750 ;
        RECT 14.555 1.580 14.725 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
        RECT 15.515 -0.085 15.685 0.085 ;
        RECT 15.995 -0.085 16.165 0.085 ;
        RECT 16.475 -0.085 16.645 0.085 ;
      LAYER met1 ;
        RECT 2.495 1.735 2.785 1.780 ;
        RECT 14.495 1.735 14.785 1.780 ;
        RECT 2.495 1.595 14.785 1.735 ;
        RECT 2.495 1.550 2.785 1.595 ;
        RECT 14.495 1.550 14.785 1.595 ;
  END
END sky130_fd_sc_hs__sedfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hs__tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hs__tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.480 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 0.455 1.275 ;
        RECT 0.000 0.000 0.480 0.245 ;
      LAYER li1 ;
        RECT 0.090 0.265 0.390 1.440 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 0.670 3.520 ;
      LAYER li1 ;
        RECT 0.090 1.890 0.390 3.065 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.480 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.480 3.415 ;
        RECT 0.000 -0.085 0.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
  END
END sky130_fd_sc_hs__tap_1

#--------EOF---------

MACRO sky130_fd_sc_hs__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hs__tap_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.960 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 0.935 1.275 ;
        RECT 0.000 0.000 0.960 0.245 ;
      LAYER li1 ;
        RECT 0.090 0.265 0.870 1.440 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.150 3.520 ;
      LAYER li1 ;
        RECT 0.090 1.890 0.870 3.065 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.960 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.960 3.415 ;
        RECT 0.000 -0.085 0.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
  END
END sky130_fd_sc_hs__tap_2

#--------EOF---------

MACRO sky130_fd_sc_hs__tapmet1_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hs__tapmet1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.245 0.935 1.275 ;
        RECT 0.000 0.000 0.960 0.245 ;
      LAYER met1 ;
        RECT 0.080 0.425 0.400 0.685 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 0.960 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 1.150 3.520 ;
      LAYER met1 ;
        RECT 0.560 2.645 0.880 2.905 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.960 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.960 3.415 ;
        RECT 0.090 2.210 0.870 3.065 ;
        RECT 0.090 0.265 0.870 1.105 ;
        RECT 0.000 -0.085 0.960 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 0.635 2.690 0.805 2.860 ;
        RECT 0.155 0.470 0.325 0.640 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
  END
END sky130_fd_sc_hs__tapmet1_2

#--------EOF---------

MACRO sky130_fd_sc_hs__tapvgnd2_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hs__tapvgnd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.190 0.455 1.275 ;
      LAYER met1 ;
        RECT 0.000 -0.245 0.480 0.245 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 0.670 3.520 ;
      LAYER met1 ;
        RECT 0.080 2.275 0.400 2.535 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.480 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.480 3.415 ;
        RECT 0.090 1.890 0.390 3.065 ;
        RECT 0.090 0.085 0.390 1.440 ;
        RECT 0.000 -0.085 0.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.155 2.320 0.325 2.490 ;
        RECT 0.155 -0.085 0.325 0.085 ;
  END
END sky130_fd_sc_hs__tapvgnd2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__tapvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hs__tapvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.190 0.455 1.275 ;
      LAYER met1 ;
        RECT 0.000 -0.245 0.480 0.245 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 0.670 3.520 ;
      LAYER met1 ;
        RECT 0.080 2.645 0.400 2.905 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 0.480 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.480 3.415 ;
        RECT 0.090 1.890 0.390 3.065 ;
        RECT 0.090 0.085 0.390 1.440 ;
        RECT 0.000 -0.085 0.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.155 2.690 0.325 2.860 ;
        RECT 0.155 -0.085 0.325 0.085 ;
  END
END sky130_fd_sc_hs__tapvgnd_1

#--------EOF---------

MACRO sky130_fd_sc_hs__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hs__tapvpwrvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.480 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.190 0.455 1.275 ;
      LAYER met1 ;
        RECT 0.000 -0.245 0.480 0.245 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 0.670 3.520 ;
      LAYER met1 ;
        RECT 0.000 3.085 0.480 3.575 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 0.480 3.415 ;
        RECT 0.090 2.205 0.390 3.245 ;
        RECT 0.090 0.085 0.390 1.105 ;
        RECT 0.000 -0.085 0.480 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
  END
END sky130_fd_sc_hs__tapvpwrvgnd_1

#--------EOF---------

MACRO sky130_fd_sc_hs__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.350 1.845 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.501000 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.950 2.185 2.120 ;
        RECT 1.175 1.780 1.345 1.950 ;
        RECT 0.945 1.435 1.345 1.780 ;
        RECT 2.015 1.680 2.185 1.950 ;
        RECT 2.015 1.350 2.465 1.680 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.360 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 1.325 1.365 ;
        RECT 0.005 0.245 3.335 1.240 ;
        RECT 0.000 0.000 3.360 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 3.550 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.360 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.699800 ;
    PORT
      LAYER li1 ;
        RECT 2.045 2.290 2.685 2.980 ;
        RECT 2.355 2.020 2.685 2.290 ;
        RECT 2.355 1.850 3.275 2.020 ;
        RECT 3.105 1.130 3.275 1.850 ;
        RECT 2.975 0.350 3.275 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.360 3.415 ;
        RECT 0.175 2.290 0.505 3.245 ;
        RECT 0.175 1.905 0.425 2.290 ;
        RECT 0.675 2.120 1.005 2.785 ;
        RECT 1.415 2.290 1.745 3.245 ;
        RECT 2.855 2.190 3.185 3.245 ;
        RECT 0.605 1.950 1.005 2.120 ;
        RECT 0.605 1.255 0.775 1.950 ;
        RECT 2.635 1.300 2.935 1.630 ;
        RECT 0.105 0.085 0.435 1.255 ;
        RECT 0.605 1.180 1.225 1.255 ;
        RECT 2.635 1.180 2.805 1.300 ;
        RECT 0.605 1.085 2.805 1.180 ;
        RECT 0.895 1.010 2.805 1.085 ;
        RECT 0.895 0.575 1.225 1.010 ;
        RECT 1.435 0.670 2.770 0.840 ;
        RECT 1.435 0.510 1.765 0.670 ;
        RECT 2.440 0.510 2.770 0.670 ;
        RECT 1.935 0.085 2.265 0.500 ;
        RECT 0.000 -0.085 3.360 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
  END
END sky130_fd_sc_hs__xnor2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.819000 ;
    PORT
      LAYER met1 ;
        RECT 0.575 1.365 0.865 1.410 ;
        RECT 2.975 1.365 3.265 1.410 ;
        RECT 0.575 1.225 3.265 1.365 ;
        RECT 0.575 1.180 0.865 1.225 ;
        RECT 2.975 1.180 3.265 1.225 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.819000 ;
    PORT
      LAYER li1 ;
        RECT 2.605 2.060 5.195 2.230 ;
        RECT 2.605 1.890 2.775 2.060 ;
        RECT 1.345 1.720 2.775 1.890 ;
        RECT 1.345 1.350 1.675 1.720 ;
        RECT 3.925 1.180 4.255 1.550 ;
        RECT 5.025 1.180 5.195 2.060 ;
        RECT 3.925 1.010 5.195 1.180 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 5.280 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.225 1.030 5.240 1.240 ;
        RECT 0.225 0.780 5.275 1.030 ;
        RECT 0.005 0.245 5.275 0.780 ;
        RECT 0.000 0.000 5.280 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 5.470 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 5.280 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.072800 ;
    PORT
      LAYER li1 ;
        RECT 2.045 2.570 2.435 2.980 ;
        RECT 3.805 2.570 4.135 2.735 ;
        RECT 2.045 2.490 4.135 2.570 ;
        RECT 0.085 2.400 4.135 2.490 ;
        RECT 0.085 2.320 2.435 2.400 ;
        RECT 0.085 1.010 0.255 2.320 ;
        RECT 2.045 2.060 2.435 2.320 ;
        RECT 0.085 0.840 0.835 1.010 ;
        RECT 0.665 0.425 0.835 0.840 ;
        RECT 2.190 0.425 2.575 0.500 ;
        RECT 0.665 0.255 2.575 0.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 5.280 3.415 ;
        RECT 0.115 2.660 0.445 3.245 ;
        RECT 1.230 2.660 1.875 3.245 ;
        RECT 2.640 2.740 2.970 3.245 ;
        RECT 3.260 2.905 4.635 3.075 ;
        RECT 3.260 2.740 3.600 2.905 ;
        RECT 4.305 2.400 4.635 2.905 ;
        RECT 4.805 2.400 5.135 3.245 ;
        RECT 0.650 1.820 1.175 2.150 ;
        RECT 0.425 1.180 0.835 1.550 ;
        RECT 1.005 1.180 1.175 1.820 ;
        RECT 3.025 1.720 4.675 1.890 ;
        RECT 3.025 1.550 3.355 1.720 ;
        RECT 1.915 1.180 2.585 1.550 ;
        RECT 3.005 1.180 3.355 1.550 ;
        RECT 4.445 1.680 4.675 1.720 ;
        RECT 4.445 1.350 4.855 1.680 ;
        RECT 1.005 1.010 2.585 1.180 ;
        RECT 0.115 0.085 0.495 0.670 ;
        RECT 1.005 0.635 1.450 1.010 ;
        RECT 2.755 0.840 3.085 1.010 ;
        RECT 1.680 0.670 5.165 0.840 ;
        RECT 1.680 0.595 2.010 0.670 ;
        RECT 2.755 0.350 3.085 0.670 ;
        RECT 3.265 0.085 3.600 0.500 ;
        RECT 3.780 0.490 4.110 0.670 ;
        RECT 4.310 0.085 4.655 0.500 ;
        RECT 4.835 0.490 5.165 0.670 ;
        RECT 0.000 -0.085 5.280 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 0.635 1.210 0.805 1.380 ;
        RECT 3.035 1.210 3.205 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
  END
END sky130_fd_sc_hs__xnor2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.735 1.345 1.780 ;
        RECT 4.415 1.735 4.705 1.780 ;
        RECT 1.055 1.595 4.705 1.735 ;
        RECT 1.055 1.550 1.345 1.595 ;
        RECT 4.415 1.550 4.705 1.595 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.945 6.535 2.115 ;
        RECT 1.985 1.680 2.155 1.945 ;
        RECT 1.485 1.350 2.155 1.680 ;
        RECT 6.365 1.765 6.535 1.945 ;
        RECT 6.365 1.350 8.155 1.765 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.425 1.140 9.115 1.240 ;
        RECT 0.005 0.245 9.115 1.140 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.474200 ;
    PORT
      LAYER li1 ;
        RECT 7.325 2.455 7.655 2.735 ;
        RECT 2.545 2.285 7.655 2.455 ;
        RECT 7.325 2.105 7.655 2.285 ;
        RECT 8.225 2.105 8.555 2.735 ;
        RECT 7.325 1.935 8.555 2.105 ;
        RECT 8.325 1.180 8.495 1.935 ;
        RECT 3.035 1.010 8.495 1.180 ;
        RECT 3.035 0.595 3.365 1.010 ;
        RECT 4.060 0.595 4.390 1.010 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.115 1.820 0.365 3.245 ;
        RECT 0.565 2.120 0.895 2.700 ;
        RECT 1.095 2.290 1.265 3.245 ;
        RECT 2.000 2.965 2.340 3.245 ;
        RECT 3.080 2.965 3.410 3.245 ;
        RECT 3.580 2.795 4.590 2.955 ;
        RECT 1.465 2.625 4.590 2.795 ;
        RECT 4.810 2.795 5.060 2.980 ;
        RECT 5.265 2.965 5.600 3.245 ;
        RECT 5.805 2.795 6.135 2.980 ;
        RECT 6.340 2.965 6.670 3.245 ;
        RECT 6.875 2.905 9.005 3.075 ;
        RECT 6.875 2.795 7.125 2.905 ;
        RECT 4.810 2.625 7.125 2.795 ;
        RECT 1.465 2.120 1.795 2.625 ;
        RECT 7.855 2.275 8.025 2.905 ;
        RECT 0.565 1.950 1.795 2.120 ;
        RECT 0.565 1.820 0.895 1.950 ;
        RECT 8.755 1.935 9.005 2.905 ;
        RECT 1.085 1.650 1.315 1.780 ;
        RECT 0.545 1.320 1.315 1.650 ;
        RECT 2.395 1.350 4.085 1.680 ;
        RECT 4.445 1.350 5.835 1.775 ;
        RECT 2.395 1.180 2.565 1.350 ;
        RECT 0.115 0.980 1.375 1.150 ;
        RECT 0.115 0.350 0.365 0.980 ;
        RECT 0.545 0.085 0.875 0.810 ;
        RECT 1.045 0.600 1.375 0.980 ;
        RECT 1.545 1.010 2.565 1.180 ;
        RECT 1.545 0.770 1.875 1.010 ;
        RECT 8.675 0.840 9.005 1.130 ;
        RECT 1.045 0.350 2.305 0.600 ;
        RECT 2.535 0.425 2.865 0.840 ;
        RECT 3.535 0.425 3.865 0.840 ;
        RECT 4.560 0.670 9.005 0.840 ;
        RECT 4.560 0.425 4.890 0.670 ;
        RECT 2.535 0.255 4.890 0.425 ;
        RECT 5.070 0.085 5.400 0.500 ;
        RECT 5.580 0.350 5.910 0.670 ;
        RECT 6.090 0.085 6.420 0.500 ;
        RECT 6.600 0.350 6.930 0.670 ;
        RECT 7.110 0.085 7.475 0.500 ;
        RECT 7.655 0.350 7.985 0.670 ;
        RECT 8.165 0.085 8.495 0.500 ;
        RECT 8.675 0.350 9.005 0.670 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 1.115 1.580 1.285 1.750 ;
        RECT 4.475 1.580 4.645 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
  END
END sky130_fd_sc_hs__xnor2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.425 7.205 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.693000 ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.350 4.375 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.350 1.325 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.160 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.355 1.370 8.155 1.375 ;
        RECT 0.005 1.140 1.665 1.360 ;
        RECT 3.285 1.140 8.155 1.370 ;
        RECT 0.005 0.245 8.155 1.140 ;
        RECT 0.000 0.000 8.160 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.350 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.160 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.530100 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.840 0.355 2.980 ;
        RECT 0.085 1.170 0.255 1.840 ;
        RECT 0.085 0.440 0.445 1.170 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.160 3.415 ;
        RECT 0.555 2.290 0.805 3.245 ;
        RECT 0.975 2.905 2.655 3.075 ;
        RECT 0.975 2.120 1.145 2.905 ;
        RECT 1.875 2.540 2.125 2.735 ;
        RECT 2.325 2.710 2.655 2.905 ;
        RECT 3.395 2.710 3.725 3.245 ;
        RECT 4.490 2.905 7.090 3.075 ;
        RECT 4.490 2.710 4.820 2.905 ;
        RECT 5.015 2.540 5.265 2.575 ;
        RECT 0.615 1.950 1.145 2.120 ;
        RECT 1.315 1.950 1.665 2.500 ;
        RECT 1.875 2.370 5.265 2.540 ;
        RECT 1.875 1.950 2.125 2.370 ;
        RECT 2.850 2.030 3.185 2.200 ;
        RECT 0.615 1.670 0.785 1.950 ;
        RECT 0.425 1.340 0.785 1.670 ;
        RECT 0.615 0.830 0.785 1.340 ;
        RECT 1.495 1.750 1.665 1.950 ;
        RECT 2.515 1.750 2.845 1.810 ;
        RECT 1.495 1.580 2.845 1.750 ;
        RECT 1.495 1.170 1.665 1.580 ;
        RECT 2.515 1.480 2.845 1.580 ;
        RECT 1.135 1.000 1.665 1.170 ;
        RECT 1.835 1.310 2.275 1.410 ;
        RECT 3.015 1.310 3.185 2.030 ;
        RECT 1.835 1.140 3.185 1.310 ;
        RECT 0.615 0.660 1.665 0.830 ;
        RECT 0.625 0.085 0.955 0.490 ;
        RECT 1.495 0.425 1.665 0.660 ;
        RECT 1.835 0.595 2.165 1.140 ;
        RECT 3.355 0.970 3.525 2.370 ;
        RECT 3.920 1.950 4.715 2.200 ;
        RECT 4.545 1.685 4.715 1.950 ;
        RECT 5.015 1.855 5.265 2.370 ;
        RECT 5.550 2.565 6.590 2.735 ;
        RECT 5.550 2.105 5.880 2.565 ;
        RECT 6.080 1.935 6.250 2.395 ;
        RECT 5.435 1.765 6.250 1.935 ;
        RECT 4.545 1.355 5.045 1.685 ;
        RECT 5.435 1.410 5.605 1.765 ;
        RECT 6.420 1.595 6.590 2.565 ;
        RECT 6.760 2.120 7.090 2.905 ;
        RECT 7.260 2.290 7.590 3.245 ;
        RECT 7.790 2.190 8.075 2.930 ;
        RECT 6.760 1.950 7.620 2.120 ;
        RECT 4.545 1.180 4.715 1.355 ;
        RECT 5.315 1.185 5.605 1.410 ;
        RECT 3.905 1.010 4.715 1.180 ;
        RECT 5.020 1.180 5.605 1.185 ;
        RECT 5.775 1.425 6.590 1.595 ;
        RECT 7.415 1.755 7.620 1.950 ;
        RECT 7.415 1.425 7.665 1.755 ;
        RECT 5.020 1.015 5.485 1.180 ;
        RECT 2.335 0.425 2.665 0.970 ;
        RECT 1.495 0.255 2.665 0.425 ;
        RECT 2.835 0.840 3.525 0.970 ;
        RECT 5.775 0.935 6.085 1.425 ;
        RECT 7.415 1.255 7.620 1.425 ;
        RECT 7.835 1.255 8.075 2.190 ;
        RECT 2.835 0.765 5.180 0.840 ;
        RECT 6.255 0.765 6.535 1.210 ;
        RECT 2.835 0.670 6.535 0.765 ;
        RECT 2.835 0.350 3.165 0.670 ;
        RECT 5.010 0.595 6.535 0.670 ;
        RECT 6.705 1.085 7.620 1.255 ;
        RECT 3.395 0.085 3.725 0.500 ;
        RECT 4.465 0.425 4.840 0.500 ;
        RECT 6.705 0.425 7.035 1.085 ;
        RECT 4.465 0.255 7.035 0.425 ;
        RECT 7.205 0.085 7.615 0.915 ;
        RECT 7.795 0.585 8.075 1.255 ;
        RECT 0.000 -0.085 8.160 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 2.075 1.210 2.245 1.380 ;
        RECT 5.435 1.210 5.605 1.380 ;
        RECT 5.915 1.210 6.085 1.380 ;
        RECT 7.835 1.210 8.005 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
      LAYER met1 ;
        RECT 2.015 1.365 2.305 1.410 ;
        RECT 5.375 1.365 5.665 1.410 ;
        RECT 2.015 1.225 5.665 1.365 ;
        RECT 2.015 1.180 2.305 1.225 ;
        RECT 5.375 1.180 5.665 1.225 ;
        RECT 5.855 1.365 6.145 1.410 ;
        RECT 7.775 1.365 8.065 1.410 ;
        RECT 5.855 1.225 8.065 1.365 ;
        RECT 5.855 1.180 6.145 1.225 ;
        RECT 7.775 1.180 8.065 1.225 ;
  END
END sky130_fd_sc_hs__xnor3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.375 1.315 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.693000 ;
    PORT
      LAYER li1 ;
        RECT 3.735 1.350 4.405 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.350 7.175 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.605 1.315 3.640 1.395 ;
        RECT 1.605 1.175 4.710 1.315 ;
        RECT 0.045 1.140 4.710 1.175 ;
        RECT 6.280 1.140 8.635 1.360 ;
        RECT 0.045 0.245 8.635 1.140 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 7.750 1.840 8.095 2.980 ;
        RECT 7.925 1.170 8.095 1.840 ;
        RECT 7.765 0.440 8.095 1.170 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.085 2.290 0.445 2.885 ;
        RECT 0.645 2.305 0.925 3.245 ;
        RECT 1.095 2.905 3.675 3.075 ;
        RECT 0.085 1.065 0.325 2.290 ;
        RECT 1.095 2.120 1.375 2.905 ;
        RECT 0.495 1.950 1.375 2.120 ;
        RECT 1.545 2.565 2.605 2.735 ;
        RECT 3.345 2.710 3.675 2.905 ;
        RECT 4.455 2.735 4.785 3.245 ;
        RECT 5.535 2.905 7.210 3.075 ;
        RECT 5.535 2.735 5.865 2.905 ;
        RECT 0.495 1.235 0.745 1.950 ;
        RECT 0.575 1.205 0.745 1.235 ;
        RECT 1.545 1.380 1.715 2.565 ;
        RECT 1.885 1.720 2.105 2.395 ;
        RECT 2.275 1.890 2.605 2.565 ;
        RECT 2.835 2.540 3.065 2.620 ;
        RECT 6.070 2.565 6.320 2.735 ;
        RECT 4.585 2.540 6.320 2.565 ;
        RECT 2.835 2.395 6.320 2.540 ;
        RECT 2.835 2.370 4.755 2.395 ;
        RECT 2.835 1.875 3.145 2.370 ;
        RECT 3.395 1.950 4.255 2.200 ;
        RECT 1.885 1.550 2.755 1.720 ;
        RECT 3.395 1.705 3.565 1.950 ;
        RECT 0.085 0.385 0.405 1.065 ;
        RECT 0.575 1.035 1.345 1.205 ;
        RECT 1.545 1.165 2.385 1.380 ;
        RECT 0.585 0.085 0.915 0.865 ;
        RECT 1.095 0.425 1.345 1.035 ;
        RECT 1.625 0.765 1.955 0.995 ;
        RECT 2.135 0.935 2.385 1.165 ;
        RECT 2.555 1.285 2.755 1.550 ;
        RECT 3.155 1.375 3.565 1.705 ;
        RECT 2.555 0.955 2.985 1.285 ;
        RECT 3.395 1.125 3.565 1.375 ;
        RECT 3.395 0.955 4.090 1.125 ;
        RECT 4.585 0.965 4.755 2.370 ;
        RECT 4.925 1.975 5.335 2.225 ;
        RECT 6.070 1.975 6.320 2.395 ;
        RECT 4.925 1.305 5.155 1.975 ;
        RECT 6.505 1.950 6.870 2.500 ;
        RECT 7.040 2.120 7.210 2.905 ;
        RECT 7.380 2.290 7.550 3.245 ;
        RECT 7.040 1.950 7.580 2.120 ;
        RECT 6.505 1.805 6.675 1.950 ;
        RECT 5.325 1.475 6.675 1.805 ;
        RECT 4.925 1.135 6.160 1.305 ;
        RECT 4.585 0.785 5.160 0.965 ;
        RECT 2.555 0.765 5.160 0.785 ;
        RECT 1.625 0.615 5.160 0.765 ;
        RECT 1.625 0.595 2.725 0.615 ;
        RECT 3.200 0.425 3.530 0.445 ;
        RECT 1.095 0.255 3.530 0.425 ;
        RECT 4.270 0.085 4.600 0.445 ;
        RECT 4.830 0.350 5.160 0.615 ;
        RECT 5.330 0.425 5.660 0.965 ;
        RECT 5.830 0.595 6.160 1.135 ;
        RECT 6.390 1.170 6.675 1.475 ;
        RECT 7.410 1.670 7.580 1.950 ;
        RECT 8.280 1.820 8.530 3.245 ;
        RECT 7.410 1.340 7.755 1.670 ;
        RECT 7.410 1.180 7.580 1.340 ;
        RECT 6.390 1.000 6.720 1.170 ;
        RECT 6.890 1.010 7.580 1.180 ;
        RECT 6.890 0.830 7.060 1.010 ;
        RECT 6.330 0.660 7.060 0.830 ;
        RECT 6.330 0.425 6.500 0.660 ;
        RECT 7.230 0.490 7.585 0.840 ;
        RECT 5.330 0.255 6.500 0.425 ;
        RECT 6.900 0.085 7.585 0.490 ;
        RECT 8.275 0.085 8.525 1.250 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 1.210 0.325 1.380 ;
        RECT 1.595 1.210 1.765 1.380 ;
        RECT 2.555 1.210 2.725 1.380 ;
        RECT 4.955 1.210 5.125 1.380 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
      LAYER met1 ;
        RECT 0.095 1.365 0.385 1.410 ;
        RECT 1.535 1.365 1.825 1.410 ;
        RECT 0.095 1.225 1.825 1.365 ;
        RECT 0.095 1.180 0.385 1.225 ;
        RECT 1.535 1.180 1.825 1.225 ;
        RECT 2.495 1.365 2.785 1.410 ;
        RECT 4.895 1.365 5.185 1.410 ;
        RECT 2.495 1.225 5.185 1.365 ;
        RECT 2.495 1.180 2.785 1.225 ;
        RECT 4.895 1.180 5.185 1.225 ;
  END
END sky130_fd_sc_hs__xnor3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.915 1.375 1.315 1.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.693000 ;
    PORT
      LAYER li1 ;
        RECT 3.940 1.350 4.270 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 6.780 1.350 7.110 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.080 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.025 1.315 3.640 1.375 ;
        RECT 2.025 1.155 4.710 1.315 ;
        RECT 0.055 1.140 4.710 1.155 ;
        RECT 6.280 1.140 10.075 1.360 ;
        RECT 0.055 0.245 10.075 1.140 ;
        RECT 0.000 0.000 10.080 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.270 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.080 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 8.280 1.840 8.640 2.980 ;
        RECT 8.470 1.625 8.640 1.840 ;
        RECT 9.180 1.625 9.535 2.980 ;
        RECT 8.470 1.420 9.535 1.625 ;
        RECT 8.470 1.170 8.675 1.420 ;
        RECT 8.345 0.470 8.675 1.170 ;
        RECT 9.205 0.440 9.535 1.420 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.085 1.845 0.365 2.885 ;
        RECT 0.565 2.290 0.895 3.245 ;
        RECT 1.065 2.905 3.680 3.075 ;
        RECT 1.065 2.120 1.395 2.905 ;
        RECT 0.535 1.950 1.395 2.120 ;
        RECT 1.565 2.565 2.725 2.735 ;
        RECT 3.350 2.710 3.680 2.905 ;
        RECT 4.390 2.730 4.720 3.245 ;
        RECT 5.485 2.905 7.315 3.075 ;
        RECT 5.485 2.730 5.815 2.905 ;
        RECT 0.085 0.865 0.285 1.845 ;
        RECT 0.535 1.465 0.705 1.950 ;
        RECT 0.455 1.205 0.705 1.465 ;
        RECT 1.565 1.375 1.765 2.565 ;
        RECT 2.305 2.290 2.725 2.565 ;
        RECT 6.020 2.560 6.270 2.735 ;
        RECT 2.895 2.540 3.145 2.545 ;
        RECT 4.440 2.540 6.270 2.560 ;
        RECT 2.895 2.390 6.270 2.540 ;
        RECT 2.895 2.370 4.610 2.390 ;
        RECT 1.935 2.120 2.135 2.155 ;
        RECT 1.935 1.675 2.245 2.120 ;
        RECT 2.895 1.875 3.145 2.370 ;
        RECT 3.600 1.950 4.270 2.200 ;
        RECT 3.600 1.705 3.770 1.950 ;
        RECT 1.935 1.505 2.755 1.675 ;
        RECT 1.595 1.335 1.765 1.375 ;
        RECT 0.455 1.035 1.425 1.205 ;
        RECT 1.595 1.165 2.385 1.335 ;
        RECT 0.085 0.365 0.495 0.865 ;
        RECT 0.665 0.085 0.995 0.865 ;
        RECT 1.175 0.425 1.425 1.035 ;
        RECT 1.625 0.765 1.955 0.995 ;
        RECT 2.135 0.935 2.385 1.165 ;
        RECT 2.555 1.205 2.755 1.505 ;
        RECT 2.995 1.375 3.770 1.705 ;
        RECT 2.555 0.955 3.020 1.205 ;
        RECT 3.600 1.125 3.770 1.375 ;
        RECT 3.600 0.955 4.090 1.125 ;
        RECT 4.440 1.030 4.610 2.370 ;
        RECT 4.780 1.950 5.280 2.220 ;
        RECT 6.020 1.970 6.270 2.390 ;
        RECT 6.440 1.990 6.960 2.500 ;
        RECT 7.130 2.120 7.315 2.905 ;
        RECT 7.485 2.290 8.110 3.245 ;
        RECT 4.780 1.380 4.950 1.950 ;
        RECT 5.120 1.720 5.450 1.780 ;
        RECT 6.440 1.720 6.610 1.990 ;
        RECT 7.130 1.950 7.490 2.120 ;
        RECT 5.120 1.550 6.610 1.720 ;
        RECT 4.780 1.210 6.160 1.380 ;
        RECT 5.405 1.180 6.160 1.210 ;
        RECT 4.440 0.785 5.160 1.030 ;
        RECT 2.555 0.765 5.160 0.785 ;
        RECT 1.625 0.615 5.160 0.765 ;
        RECT 1.625 0.595 2.725 0.615 ;
        RECT 3.200 0.425 3.530 0.445 ;
        RECT 1.175 0.255 3.530 0.425 ;
        RECT 4.270 0.085 4.600 0.445 ;
        RECT 4.830 0.350 5.160 0.615 ;
        RECT 5.330 0.425 5.660 1.010 ;
        RECT 5.830 0.595 6.160 1.180 ;
        RECT 6.390 1.170 6.610 1.550 ;
        RECT 7.320 1.670 7.490 1.950 ;
        RECT 7.685 1.840 8.110 2.290 ;
        RECT 8.810 1.820 8.980 3.245 ;
        RECT 9.710 1.820 9.960 3.245 ;
        RECT 7.320 1.340 8.300 1.670 ;
        RECT 7.320 1.180 7.490 1.340 ;
        RECT 6.390 1.000 6.720 1.170 ;
        RECT 6.890 1.010 7.490 1.180 ;
        RECT 6.890 0.830 7.060 1.010 ;
        RECT 7.915 0.840 8.165 1.170 ;
        RECT 6.330 0.660 7.060 0.830 ;
        RECT 6.330 0.425 6.500 0.660 ;
        RECT 7.230 0.490 8.165 0.840 ;
        RECT 5.330 0.255 6.500 0.425 ;
        RECT 6.900 0.085 8.165 0.490 ;
        RECT 8.855 0.085 9.025 1.250 ;
        RECT 9.715 0.085 9.965 1.250 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 0.155 1.950 0.325 2.120 ;
        RECT 1.595 1.950 1.765 2.120 ;
        RECT 2.075 1.950 2.245 2.120 ;
        RECT 4.955 1.950 5.125 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
      LAYER met1 ;
        RECT 0.095 2.105 0.385 2.150 ;
        RECT 1.535 2.105 1.825 2.150 ;
        RECT 0.095 1.965 1.825 2.105 ;
        RECT 0.095 1.920 0.385 1.965 ;
        RECT 1.535 1.920 1.825 1.965 ;
        RECT 2.015 2.105 2.305 2.150 ;
        RECT 4.895 2.105 5.185 2.150 ;
        RECT 2.015 1.965 5.185 2.105 ;
        RECT 2.015 1.920 2.305 1.965 ;
        RECT 4.895 1.920 5.185 1.965 ;
  END
END sky130_fd_sc_hs__xnor3_4

#--------EOF---------

MACRO sky130_fd_sc_hs__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 0.775 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.695 2.845 1.780 ;
        RECT 1.285 1.365 2.845 1.695 ;
        RECT 2.515 1.350 2.845 1.365 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 3.840 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.085 0.245 3.770 1.305 ;
        RECT 0.000 0.000 3.840 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.030 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 3.840 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.697200 ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.820 3.755 2.980 ;
        RECT 3.585 1.150 3.755 1.820 ;
        RECT 2.525 0.980 3.755 1.150 ;
        RECT 2.525 0.415 2.970 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 3.840 3.415 ;
        RECT 0.325 1.940 0.655 3.245 ;
        RECT 0.945 2.120 1.525 2.980 ;
        RECT 1.755 2.460 2.085 2.980 ;
        RECT 2.255 2.650 2.695 3.245 ;
        RECT 2.865 2.460 3.195 2.980 ;
        RECT 1.755 2.290 3.195 2.460 ;
        RECT 0.945 1.950 3.195 2.120 ;
        RECT 0.945 1.040 1.115 1.950 ;
        RECT 3.025 1.650 3.195 1.950 ;
        RECT 3.025 1.320 3.415 1.650 ;
        RECT 0.175 0.085 0.775 0.990 ;
        RECT 0.945 0.710 1.640 1.040 ;
        RECT 1.820 0.085 2.150 1.195 ;
        RECT 3.210 0.085 3.540 0.745 ;
        RECT 0.000 -0.085 3.840 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END sky130_fd_sc_hs__xor2_1

#--------EOF---------

MACRO sky130_fd_sc_hs__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.804000 ;
    PORT
      LAYER li1 ;
        RECT 0.585 1.620 2.515 1.790 ;
        RECT 0.585 1.165 0.915 1.620 ;
        RECT 1.845 1.350 2.515 1.620 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.804000 ;
    PORT
      LAYER li1 ;
        RECT 1.155 1.180 1.485 1.450 ;
        RECT 3.485 1.180 4.145 1.550 ;
        RECT 1.155 1.010 4.145 1.180 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 4.800 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.465 1.140 4.795 1.240 ;
        RECT 0.005 0.245 4.795 1.140 ;
        RECT 0.000 0.000 4.800 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 4.990 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 4.800 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.754100 ;
    PORT
      LAYER li1 ;
        RECT 3.025 2.020 3.195 2.735 ;
        RECT 3.025 1.850 4.685 2.020 ;
        RECT 4.355 0.840 4.685 1.850 ;
        RECT 3.330 0.670 4.685 0.840 ;
        RECT 3.330 0.595 3.660 0.670 ;
        RECT 4.355 0.350 4.685 0.670 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 4.800 3.415 ;
        RECT 0.115 2.300 0.445 3.245 ;
        RECT 1.065 2.130 1.315 2.980 ;
        RECT 1.545 2.470 1.795 2.980 ;
        RECT 1.995 2.640 2.325 3.245 ;
        RECT 2.495 2.905 3.675 3.075 ;
        RECT 2.495 2.470 2.825 2.905 ;
        RECT 1.545 2.300 2.825 2.470 ;
        RECT 3.395 2.360 3.675 2.905 ;
        RECT 3.845 2.530 4.175 3.245 ;
        RECT 4.345 2.360 4.685 2.980 ;
        RECT 3.395 2.190 4.685 2.360 ;
        RECT 0.245 1.960 2.855 2.130 ;
        RECT 0.245 0.840 0.415 1.960 ;
        RECT 2.685 1.680 2.855 1.960 ;
        RECT 2.685 1.350 3.125 1.680 ;
        RECT 0.245 0.670 1.220 0.840 ;
        RECT 0.115 0.085 0.710 0.500 ;
        RECT 0.890 0.350 1.220 0.670 ;
        RECT 1.390 0.085 1.720 0.840 ;
        RECT 1.970 0.670 3.160 0.840 ;
        RECT 1.970 0.350 2.300 0.670 ;
        RECT 2.480 0.085 2.820 0.500 ;
        RECT 2.990 0.425 3.160 0.670 ;
        RECT 3.840 0.425 4.175 0.500 ;
        RECT 2.990 0.255 4.175 0.425 ;
        RECT 0.000 -0.085 4.800 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
  END
END sky130_fd_sc_hs__xor2_2

#--------EOF---------

MACRO sky130_fd_sc_hs__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.638000 ;
    PORT
      LAYER li1 ;
        RECT 0.440 1.420 1.110 1.750 ;
        RECT 3.965 1.520 5.635 1.775 ;
        RECT 0.515 0.750 0.685 1.420 ;
        RECT 3.765 1.350 5.635 1.520 ;
        RECT 3.765 1.190 3.935 1.350 ;
        RECT 2.870 1.020 3.935 1.190 ;
        RECT 2.870 0.770 3.040 1.020 ;
        RECT 1.275 0.750 3.040 0.770 ;
        RECT 0.515 0.600 3.040 0.750 ;
        RECT 0.515 0.580 1.445 0.600 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.638000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 2.020 5.975 2.115 ;
        RECT 2.030 1.945 5.975 2.020 ;
        RECT 2.030 1.850 3.655 1.945 ;
        RECT 2.030 1.470 2.360 1.850 ;
        RECT 5.805 1.780 5.975 1.945 ;
        RECT 5.805 1.550 8.165 1.780 ;
        RECT 5.885 1.350 8.165 1.550 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 8.640 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.240 4.245 1.360 ;
        RECT 0.005 0.245 8.635 1.240 ;
        RECT 0.000 0.000 8.640 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 8.830 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 8.640 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.504500 ;
    PORT
      LAYER li1 ;
        RECT 2.985 2.455 3.315 2.735 ;
        RECT 3.885 2.455 4.215 2.735 ;
        RECT 2.985 2.285 6.315 2.455 ;
        RECT 2.985 2.190 3.315 2.285 ;
        RECT 6.145 2.120 6.315 2.285 ;
        RECT 6.145 1.950 8.505 2.120 ;
        RECT 8.335 1.180 8.505 1.950 ;
        RECT 4.105 1.010 8.505 1.180 ;
        RECT 4.105 0.850 4.275 1.010 ;
        RECT 3.210 0.680 4.275 0.850 ;
        RECT 3.210 0.470 3.540 0.680 ;
        RECT 6.835 0.595 7.165 1.010 ;
        RECT 7.845 0.595 8.015 1.010 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 8.640 3.415 ;
        RECT 0.160 2.090 0.490 2.980 ;
        RECT 0.690 2.260 0.940 3.245 ;
        RECT 1.110 2.905 2.340 3.075 ;
        RECT 1.110 2.090 1.360 2.905 ;
        RECT 0.160 1.920 1.360 2.090 ;
        RECT 0.095 0.085 0.345 1.250 ;
        RECT 0.855 1.190 1.105 1.250 ;
        RECT 1.560 1.190 1.810 2.735 ;
        RECT 2.010 2.190 2.340 2.905 ;
        RECT 2.535 2.905 4.665 3.075 ;
        RECT 4.855 2.965 5.185 3.245 ;
        RECT 2.535 2.190 2.785 2.905 ;
        RECT 3.515 2.625 3.685 2.905 ;
        RECT 4.415 2.795 4.665 2.905 ;
        RECT 5.375 2.795 5.705 2.980 ;
        RECT 5.890 2.965 6.220 3.245 ;
        RECT 6.485 2.795 6.655 2.980 ;
        RECT 4.415 2.625 6.655 2.795 ;
        RECT 6.855 2.630 7.105 3.245 ;
        RECT 6.485 2.460 6.655 2.625 ;
        RECT 7.305 2.460 7.635 2.980 ;
        RECT 7.835 2.630 8.005 3.245 ;
        RECT 8.205 2.460 8.535 2.980 ;
        RECT 6.485 2.290 8.535 2.460 ;
        RECT 2.530 1.360 3.595 1.680 ;
        RECT 2.530 1.190 2.700 1.360 ;
        RECT 0.855 0.940 2.700 1.190 ;
        RECT 0.855 0.920 1.105 0.940 ;
        RECT 4.445 0.670 6.655 0.840 ;
        RECT 1.285 0.085 1.615 0.410 ;
        RECT 2.415 0.085 2.745 0.430 ;
        RECT 3.720 0.085 4.135 0.510 ;
        RECT 4.445 0.350 4.695 0.670 ;
        RECT 4.875 0.085 5.205 0.500 ;
        RECT 5.385 0.350 5.715 0.670 ;
        RECT 5.895 0.085 6.225 0.500 ;
        RECT 6.405 0.425 6.655 0.670 ;
        RECT 7.335 0.425 7.665 0.840 ;
        RECT 8.195 0.425 8.525 0.840 ;
        RECT 6.405 0.255 8.525 0.425 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
  END
END sky130_fd_sc_hs__xor2_4

#--------EOF---------

MACRO sky130_fd_sc_hs__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.120 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.960 1.180 1.285 1.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.693000 ;
    PORT
      LAYER li1 ;
        RECT 4.920 1.350 5.250 1.780 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 6.875 1.180 7.205 1.685 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.120 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.200 1.815 1.440 ;
        RECT 3.195 1.240 4.415 1.395 ;
        RECT 5.675 1.290 7.415 1.375 ;
        RECT 5.675 1.240 9.115 1.290 ;
        RECT 3.195 1.200 9.115 1.240 ;
        RECT 0.005 0.245 9.115 1.200 ;
        RECT 0.000 0.000 9.120 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.310 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.120 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER li1 ;
        RECT 8.755 0.400 9.005 2.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.120 3.415 ;
        RECT 0.085 2.260 0.600 2.980 ;
        RECT 0.770 2.260 1.100 3.245 ;
        RECT 1.370 2.905 3.895 3.075 ;
        RECT 0.085 1.300 0.255 2.260 ;
        RECT 1.370 2.090 1.700 2.905 ;
        RECT 3.725 2.755 3.895 2.905 ;
        RECT 0.425 1.940 1.700 2.090 ;
        RECT 1.930 2.565 3.555 2.735 ;
        RECT 1.930 1.940 2.260 2.565 ;
        RECT 0.425 1.920 1.625 1.940 ;
        RECT 0.425 1.470 0.750 1.920 ;
        RECT 0.085 0.830 0.445 1.300 ;
        RECT 1.455 1.000 1.625 1.920 ;
        RECT 2.430 1.430 2.760 2.395 ;
        RECT 2.965 1.875 3.215 2.395 ;
        RECT 1.795 1.260 2.760 1.430 ;
        RECT 1.795 0.830 1.965 1.260 ;
        RECT 2.590 1.090 2.760 1.260 ;
        RECT 0.085 0.660 1.965 0.830 ;
        RECT 0.085 0.650 0.445 0.660 ;
        RECT 0.625 0.085 1.195 0.490 ;
        RECT 2.135 0.460 2.385 1.090 ;
        RECT 2.590 0.630 2.850 1.090 ;
        RECT 3.020 0.460 3.215 1.875 ;
        RECT 2.135 0.290 3.215 0.460 ;
        RECT 3.385 0.425 3.555 2.565 ;
        RECT 3.725 1.905 4.395 2.755 ;
        RECT 3.725 1.435 4.055 1.735 ;
        RECT 3.725 0.765 3.895 1.435 ;
        RECT 4.225 1.265 4.395 1.905 ;
        RECT 4.065 0.935 4.395 1.265 ;
        RECT 4.580 1.130 4.750 2.980 ;
        RECT 4.950 1.950 5.200 3.245 ;
        RECT 6.025 2.905 7.605 3.075 ;
        RECT 5.405 1.990 5.855 2.840 ;
        RECT 5.405 1.950 5.625 1.990 ;
        RECT 5.420 1.360 5.625 1.950 ;
        RECT 6.025 1.820 6.195 2.905 ;
        RECT 5.805 1.530 6.195 1.820 ;
        RECT 6.365 1.550 6.705 2.735 ;
        RECT 6.875 2.025 7.205 2.735 ;
        RECT 7.435 2.525 7.605 2.905 ;
        RECT 7.435 2.195 7.985 2.525 ;
        RECT 6.875 1.855 7.645 2.025 ;
        RECT 5.420 1.190 6.365 1.360 ;
        RECT 4.580 0.765 4.805 1.130 ;
        RECT 3.725 0.595 4.805 0.765 ;
        RECT 4.975 0.850 6.025 1.020 ;
        RECT 4.975 0.425 5.145 0.850 ;
        RECT 3.385 0.255 5.145 0.425 ;
        RECT 5.315 0.085 5.565 0.680 ;
        RECT 5.775 0.425 6.025 0.850 ;
        RECT 6.195 0.765 6.365 1.190 ;
        RECT 6.535 0.935 6.705 1.550 ;
        RECT 6.885 0.765 7.305 0.925 ;
        RECT 6.195 0.595 7.305 0.765 ;
        RECT 7.475 0.425 7.645 1.855 ;
        RECT 5.775 0.255 7.645 0.425 ;
        RECT 7.815 0.860 7.985 2.195 ;
        RECT 8.225 1.950 8.555 3.245 ;
        RECT 8.255 1.350 8.585 1.780 ;
        RECT 7.815 0.400 8.065 0.860 ;
        RECT 8.245 0.085 8.575 1.180 ;
        RECT 0.000 -0.085 9.120 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 3.035 1.580 3.205 1.750 ;
        RECT 5.435 1.580 5.605 1.750 ;
        RECT 6.395 1.580 6.565 1.750 ;
        RECT 8.315 1.580 8.485 1.750 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
      LAYER met1 ;
        RECT 2.975 1.735 3.265 1.780 ;
        RECT 5.375 1.735 5.665 1.780 ;
        RECT 2.975 1.595 5.665 1.735 ;
        RECT 2.975 1.550 3.265 1.595 ;
        RECT 5.375 1.550 5.665 1.595 ;
        RECT 6.335 1.735 6.625 1.780 ;
        RECT 8.255 1.735 8.545 1.780 ;
        RECT 6.335 1.595 8.545 1.735 ;
        RECT 6.335 1.550 6.625 1.595 ;
        RECT 8.255 1.550 8.545 1.595 ;
  END
END sky130_fd_sc_hs__xor3_1

#--------EOF---------

MACRO sky130_fd_sc_hs__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.180 1.285 1.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.693000 ;
    PORT
      LAYER li1 ;
        RECT 4.920 1.180 5.250 1.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 6.875 1.180 7.125 1.685 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 9.600 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.335 1.815 1.440 ;
        RECT 3.195 1.335 4.415 1.395 ;
        RECT 0.005 1.240 4.415 1.335 ;
        RECT 6.345 1.305 7.375 1.375 ;
        RECT 5.675 1.260 7.375 1.305 ;
        RECT 5.675 1.240 9.575 1.260 ;
        RECT 0.005 0.245 9.575 1.240 ;
        RECT 0.000 0.000 9.600 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 9.790 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 9.600 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.543200 ;
    PORT
      LAYER li1 ;
        RECT 8.705 0.370 9.035 2.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 9.600 3.415 ;
        RECT 0.085 2.260 0.595 2.955 ;
        RECT 0.765 2.260 1.095 3.245 ;
        RECT 1.310 2.905 3.895 3.075 ;
        RECT 0.085 1.275 0.255 2.260 ;
        RECT 1.310 2.090 1.640 2.905 ;
        RECT 3.725 2.755 3.895 2.905 ;
        RECT 0.425 2.075 1.640 2.090 ;
        RECT 1.850 2.565 3.555 2.735 ;
        RECT 1.850 2.075 2.180 2.565 ;
        RECT 0.425 1.920 1.625 2.075 ;
        RECT 0.425 1.445 0.745 1.920 ;
        RECT 0.085 0.830 0.445 1.275 ;
        RECT 1.455 1.000 1.625 1.920 ;
        RECT 2.350 1.565 2.680 2.395 ;
        RECT 2.885 1.875 3.215 2.395 ;
        RECT 1.795 1.395 2.680 1.565 ;
        RECT 1.795 0.830 1.965 1.395 ;
        RECT 2.510 1.225 2.680 1.395 ;
        RECT 0.085 0.660 1.965 0.830 ;
        RECT 0.085 0.650 0.445 0.660 ;
        RECT 2.135 0.595 2.305 1.225 ;
        RECT 2.510 0.765 2.875 1.225 ;
        RECT 3.045 0.595 3.215 1.875 ;
        RECT 0.625 0.085 1.195 0.490 ;
        RECT 2.135 0.425 3.215 0.595 ;
        RECT 3.385 0.425 3.555 2.565 ;
        RECT 3.725 1.905 4.395 2.755 ;
        RECT 3.725 1.435 4.055 1.735 ;
        RECT 3.725 0.765 3.895 1.435 ;
        RECT 4.225 1.265 4.395 1.905 ;
        RECT 4.065 0.935 4.395 1.265 ;
        RECT 4.580 1.010 4.750 2.980 ;
        RECT 4.950 1.820 5.200 3.245 ;
        RECT 5.405 1.920 5.840 2.980 ;
        RECT 6.010 2.905 7.450 3.075 ;
        RECT 5.510 1.185 5.680 1.920 ;
        RECT 6.010 1.685 6.180 2.905 ;
        RECT 5.850 1.355 6.180 1.685 ;
        RECT 6.350 1.525 6.600 2.700 ;
        RECT 6.785 2.025 7.050 2.690 ;
        RECT 7.280 2.500 7.450 2.905 ;
        RECT 7.280 2.195 7.805 2.500 ;
        RECT 6.785 1.855 7.465 2.025 ;
        RECT 6.350 1.355 6.705 1.525 ;
        RECT 5.510 1.015 6.365 1.185 ;
        RECT 4.580 0.765 4.805 1.010 ;
        RECT 3.725 0.595 4.805 0.765 ;
        RECT 4.975 0.675 6.025 0.845 ;
        RECT 4.975 0.425 5.145 0.675 ;
        RECT 3.385 0.255 5.145 0.425 ;
        RECT 5.315 0.085 5.565 0.505 ;
        RECT 5.775 0.425 6.025 0.675 ;
        RECT 6.195 0.765 6.365 1.015 ;
        RECT 6.535 0.935 6.705 1.355 ;
        RECT 7.295 1.265 7.465 1.855 ;
        RECT 7.635 1.605 7.805 2.195 ;
        RECT 7.975 2.320 8.530 3.245 ;
        RECT 7.975 1.820 8.145 2.320 ;
        RECT 8.315 1.650 8.525 2.150 ;
        RECT 9.235 1.820 9.485 3.245 ;
        RECT 7.635 1.435 8.025 1.605 ;
        RECT 7.295 1.095 7.605 1.265 ;
        RECT 6.885 0.765 7.265 0.925 ;
        RECT 6.195 0.595 7.265 0.765 ;
        RECT 7.435 0.425 7.605 1.095 ;
        RECT 5.775 0.255 7.605 0.425 ;
        RECT 7.775 0.370 8.025 1.435 ;
        RECT 8.195 1.320 8.525 1.650 ;
        RECT 8.205 0.085 8.535 1.150 ;
        RECT 9.215 0.085 9.465 1.150 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 3.035 1.950 3.205 2.120 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 6.395 1.950 6.565 2.120 ;
        RECT 8.315 1.950 8.485 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
      LAYER met1 ;
        RECT 2.975 2.105 3.265 2.150 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 2.975 1.965 5.665 2.105 ;
        RECT 2.975 1.920 3.265 1.965 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 6.335 2.105 6.625 2.150 ;
        RECT 8.255 2.105 8.545 2.150 ;
        RECT 6.335 1.965 8.545 2.105 ;
        RECT 6.335 1.920 6.625 1.965 ;
        RECT 8.255 1.920 8.545 1.965 ;
  END
END sky130_fd_sc_hs__xor3_2

#--------EOF---------

MACRO sky130_fd_sc_hs__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.910 1.180 1.285 1.670 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.693000 ;
    PORT
      LAYER li1 ;
        RECT 4.910 1.180 5.240 1.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 6.810 1.450 7.070 1.780 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.245 10.560 0.245 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.125 1.360 4.345 1.395 ;
        RECT 0.005 1.240 4.345 1.360 ;
        RECT 5.610 1.240 7.260 1.385 ;
        RECT 0.005 0.920 7.260 1.240 ;
        RECT 8.220 0.920 10.555 1.240 ;
        RECT 0.005 0.245 10.555 0.920 ;
        RECT 0.000 0.000 10.560 0.245 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.660 10.750 3.520 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.085 10.560 3.575 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.086400 ;
    PORT
      LAYER li1 ;
        RECT 8.685 1.820 9.125 2.980 ;
        RECT 8.955 1.470 9.125 1.820 ;
        RECT 9.665 1.550 9.995 2.980 ;
        RECT 9.665 1.470 9.940 1.550 ;
        RECT 8.955 1.300 9.940 1.470 ;
        RECT 8.955 1.085 9.160 1.300 ;
        RECT 8.830 0.350 9.160 1.085 ;
        RECT 9.690 0.350 9.940 1.300 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.245 10.560 3.415 ;
        RECT 0.085 2.180 0.365 2.980 ;
        RECT 0.565 2.180 0.895 3.245 ;
        RECT 1.065 2.905 3.825 3.075 ;
        RECT 0.085 1.250 0.255 2.180 ;
        RECT 1.065 2.010 1.395 2.905 ;
        RECT 3.655 2.755 3.825 2.905 ;
        RECT 1.600 2.565 3.485 2.735 ;
        RECT 1.600 2.180 1.930 2.565 ;
        RECT 0.425 1.840 1.625 2.010 ;
        RECT 0.425 1.470 0.700 1.840 ;
        RECT 0.085 0.750 0.445 1.250 ;
        RECT 1.455 0.920 1.625 1.840 ;
        RECT 2.135 1.590 2.385 2.395 ;
        RECT 2.555 1.875 3.145 2.395 ;
        RECT 1.795 1.420 2.805 1.590 ;
        RECT 1.795 0.750 1.965 1.420 ;
        RECT 0.085 0.580 1.965 0.750 ;
        RECT 2.135 0.620 2.385 1.250 ;
        RECT 2.555 0.790 2.805 1.420 ;
        RECT 2.975 0.620 3.145 1.875 ;
        RECT 0.085 0.570 0.445 0.580 ;
        RECT 2.135 0.450 3.145 0.620 ;
        RECT 3.315 0.425 3.485 2.565 ;
        RECT 3.655 1.905 4.325 2.755 ;
        RECT 3.655 1.435 3.985 1.735 ;
        RECT 3.655 0.765 3.825 1.435 ;
        RECT 4.155 1.265 4.325 1.905 ;
        RECT 3.995 0.935 4.325 1.265 ;
        RECT 4.535 1.130 4.705 2.980 ;
        RECT 4.905 1.820 5.235 3.245 ;
        RECT 5.965 2.905 7.500 3.075 ;
        RECT 5.405 1.920 5.795 2.800 ;
        RECT 5.435 1.290 5.605 1.920 ;
        RECT 5.965 1.750 6.135 2.905 ;
        RECT 6.305 1.920 6.640 2.735 ;
        RECT 6.835 2.120 7.085 2.735 ;
        RECT 7.330 2.710 7.500 2.905 ;
        RECT 7.330 2.290 7.750 2.710 ;
        RECT 6.835 1.950 7.410 2.120 ;
        RECT 5.775 1.460 6.135 1.750 ;
        RECT 4.535 0.765 4.740 1.130 ;
        RECT 5.435 1.120 6.300 1.290 ;
        RECT 3.655 0.595 4.740 0.765 ;
        RECT 4.910 0.780 5.960 0.950 ;
        RECT 4.910 0.425 5.080 0.780 ;
        RECT 0.625 0.085 1.035 0.410 ;
        RECT 3.315 0.255 5.080 0.425 ;
        RECT 5.250 0.085 5.500 0.610 ;
        RECT 5.710 0.425 5.960 0.780 ;
        RECT 6.130 0.765 6.300 1.120 ;
        RECT 6.470 0.935 6.640 1.920 ;
        RECT 6.820 0.765 7.070 1.275 ;
        RECT 6.130 0.595 7.070 0.765 ;
        RECT 7.240 0.425 7.410 1.950 ;
        RECT 5.710 0.255 7.410 0.425 ;
        RECT 7.580 0.745 7.750 2.290 ;
        RECT 7.945 2.330 8.500 3.245 ;
        RECT 7.945 1.820 8.115 2.330 ;
        RECT 8.285 1.585 8.515 2.150 ;
        RECT 9.295 1.820 9.465 3.245 ;
        RECT 10.195 1.820 10.445 3.245 ;
        RECT 7.920 1.255 8.785 1.585 ;
        RECT 7.580 0.415 8.150 0.745 ;
        RECT 8.330 0.085 8.660 1.085 ;
        RECT 9.340 0.085 9.510 1.130 ;
        RECT 10.120 0.085 10.450 1.130 ;
        RECT 0.000 -0.085 10.560 0.085 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 2.555 1.950 2.725 2.120 ;
        RECT 5.435 1.950 5.605 2.120 ;
        RECT 6.395 1.950 6.565 2.120 ;
        RECT 8.315 1.950 8.485 2.120 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
      LAYER met1 ;
        RECT 2.495 2.105 2.785 2.150 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 2.495 1.965 5.665 2.105 ;
        RECT 2.495 1.920 2.785 1.965 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 6.335 2.105 6.625 2.150 ;
        RECT 8.255 2.105 8.545 2.150 ;
        RECT 6.335 1.965 8.545 2.105 ;
        RECT 6.335 1.920 6.625 1.965 ;
        RECT 8.255 1.920 8.545 1.965 ;
  END
END sky130_fd_sc_hs__xor3_4

#--------EOF---------


END LIBRARY
